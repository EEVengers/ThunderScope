`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mVY97ltKYXBVEfL1P9h8p9hjEMR9ha4yGYTC4H02CeaLQS43wrYOCKyQk7quiMIb78kvKcaNj/LI
+uA+n7B67w==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
q7G86K8lWbpUfI4MpktD23vIx55ffXnFlN8f2h9XlaWqH5Qusw0/DKgmu2Eoc6b4nIdM87lvf7E+
nRLq7mHUsUt9DFqDHcv5KzjO5zVBw0HjdoowHARfuIv8Ssr+qDOCb2jFoDJoItDJZJlzpM5Jl/Or
eJDr63/KIW9EP2fsoKI=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e3zjJPnG9T9FyqIwJm/mLt2Fkj+06G1l61KBXHN6ASIUPeeaGVO9kFatWwk8pwbPK9WohVCdrR8C
W5cSIZ3EwNd7lYt1FASCBTjDeruo/1gbwXq7wMq3HtpODMdrnkrS4s/hYG7Zx2IFFQLdSy+LC+4O
zDozhIDto8mR5ORHW6LAQxOQ0rUPTAaKJzYEJkOqGSW0KidL0cIrs0CmLr3HxrJH9mIid873DgjB
+Qfs5LuHTMQ8PsOZzYiVfzyO2H367cY79HDp6G5VodHvc9xu8CTADwoEsTfJmZFTGLhXMnwqWGEc
qSR6YXiYhTwkfB+fS6W2G7Mgve3Suca2G+b8yg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LsGXMukryreLoI5Hles5lL14zMoDfWMgbDmnDJpX4Qe3LlBUO/Wh15G3gCvUZnabcxk+09Sb6wV2
H7sC+5q96wUad64SXdm1y7vO7/D4mQP8ltYzaFqUGvUpWel4xeVyFgXejA443xGnMtn/o3JRLm5g
I+pO/shphPYN1TJTcqAF/tPb7Q2E/jd2MiPmjVT+nR8K0sx9jG81DAd1OgrMpuMhAMDSw4YQLrip
5QFq3GuHotMnPfPioR7uGTZixHvhA4YeWDRPUtcz4MIwMgWgENlhmEYx259gKEHs0dCJMfOIb6kw
7OdukzaTDVRsjdq0TWuMKAmX6jL2UAx48k/yKg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bxr1j6oyTJljxhJxpMr1uRau1xfBc+cki6VAt6sMd3BAoXo3ClmSMux159539ZcL5/aK1Dr7B3QJ
D7Qp0RwAVoGHFreIXlBSZVonkUKq3+7CQ9yFby0sfH/tK39wRuaRVeSqUwnn01PUaJJpRntyBwmT
TKB6Mbj/+lwnC2yUEKg=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T8Eq6oRHtKtifWXUMklw9lgD964e3iY5cI2PBI9b9cnrPfBF26I3YbQPJF84fAZvRGtcYbrPBtuo
S/LKn09DVD+DFTtRSGcmr0xYMq7s+wRhHoMQYc8JB0nPYZxgTLNFn+3TMAo8LjQ1q0oTrXLzfL/6
kV5l2vCn5EfcFtaoUy9id3cGUqkzKqHDr115FzTg93a8xMIKzpJ2KHE6Mm7BLD6dxaoFSCSJlQiH
1Tkf7YOSdhlDUpdUaQLfyHLu8YMeWNll0eVnjdpkP+0mTrWri3gWtE3mvuoOvZwTSJ49+14SmXSg
VTmKQhEEn6tVTandnvsOXAll1/nR32q/NTQIvw==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BgFAkc/v6hlsJtYz/aYJ2DP1ljfvs1Tlg4yukDxwReed6Sw2BjGDKFVZjvXWq4BFQ0/0srmPlmzs
PEoPl7iP+/sSnD3DqDs5eKA0Ife8HRhdLVUktuVbNp+GLh6Kf/ur1HpPjxOh09G4sWsTknUF5Z45
ychiaPlvmpkDjCflUSbGdUadg1UATICEvYRQ7Ai9ZLXRcE9tIC9mJG9RAembmKsbfbPhA9pn9u6Z
+wJXU7yFsQG54IIxZA1/5RuRlhdhpia+/mzXqNLkTIGX4n92k8irzVg2rPLjhUunVETega6zdShV
60B8B5bVZkrKvlrhHa0v1xc1mKlkhplK/YRP6A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aJu+3gyuKQkNQj/ks1jmFhEdXMwCEftkOwUsy/D0XW6id51ySnG0zSvYudQgvuou0LJ8DVDTx+bL
vJDV14tuU9OpG2vIOwMhK/5hKPq6TCYb/MDNMt4vxUKDsaQmi7KHcf8AgTR+iJi1e6R8vlzURx2b
MpRDDvF78OfOi/cjxV8U8xH8QbBjEJDuMB0kw40UDxY12FxSGUkBA5X+tMBAjOQEiw9kwHw1f5He
BSyq9HXpwHqCFJUmNhs7Y5i00yY8oiVPssk9Mriko4At+1EKXPKjpdfQjCvvCxzBmF+qcEw8J0H9
gd0Zj6Cyes/d0AvHnTisyRxTxVwatFa+eqRPgg==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JaKk9Ld24oYI7V/2d1srKafZr5tqcWioYxrKT5vcL5rc4tI9DH50dLZ0ObXO5SbSg8XqVNSorfCC
QDDw05Z5Q8ll658UCz1bRjBG8cclvWRWj1FFNvsXeIJ/IhGAfa0M7q9QkYSGn1b4y2cvSCrE3GRT
iX1VWHhqjKOROe/Z1paEeTpdQ9Aak/W1J50cUqxG5ijKU6mZtpRL/r3SqwsXTq2bY6CNbPqLrELS
4O86bIke4tv/TTnqntgxNrWgtjG7aCLkrGLGHuJf/YzR5UqkgLlzCWFLEbHteHxqNkMeYRCEWjTN
EOxEY5E2QmnyBAGLHEvsPhvjKcwUPeZ3oiQSOA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1069024)
`protect data_block
pslSeULstnh2ViYIoN8Yv9llrnk49XkLLRD0cNF3Ety5HblZL932QqdcpLgmT34scWEpQHxP+N1X
9xJhwc57NrKmdD4hCVOKVTnCVPXJCFdf1hnIatFFF7sTTGcTxdhspK5mrVoeQKD+AqraWvBnQfPT
624tvsSJgiOPMD9Be94YTt4PCEq5u0DUlkw/GRyoRP0eeKe1+V5813Sj99M327EECG5goizkgOfS
yVByYIbt7GP/3PN9HRXNIfgVjqC5ZVz1FhFiJNT9L/KYAes3UY2WBH9uvIqrU7mcEeK1aNckn8u+
/vM6Jzozn4ATDPVd8e1aPbGLPw22JRXqy94HVQgjzaLF01rAJaNxjwIQkaUF6PgigXx/I2FPM/m4
uMsvg/LBN7BQWwwT3IZggA37BIciMgfhVBzHFtQafzD9OOQ46EQNxdpEaACNORqEWZcdoF0xsafy
iwOvHqv6LggWIR/t/4tLD4Lr10dukSig6T4KPL+B3r8DK9jGCKrBM8jHL1WJ4j0uTSsx28dRG29M
9TM4uzsau8qHVq32ANkE9o3SbkMhio1LFMgI9vbUzXFgjsDBE/boJsJBqD9n37DVyK8aT44FsB+B
dx+vzXf1l/Pbi9Aa2iBhIxhmVbGXAwQr9EQpEhwcKDJgpjhInkp0s8loeZR4Ldwyl41jfF45UKwf
m9vjV4x/FUH9Tyef+S9HRdNof+j6O42CI44OMZJLtAGqiU/WGfhmJ9elEuwh1EGYhME8FQV6QlB+
YI4Oy+mzixXqnYByfVcbh8eteDQFOWPw18jV8RPp8s4QJBozUyBAAtDduXWsQrr+ELi1u4193d3E
RCJ5/Qh49stssDqOq0+Kq406+Zuz+75goCghSBb5O620J8s186M7i4kHnAHFOEVI5uwk7xhF+1DS
uJ/7VHgzj6YCtYM6FDXPua+aOhXGXijaI3UYXXOuziZazvDr6ZCJ8dtvj9UTKcQzl8/b7+fxjqMA
xN3H6DyNMok6h7mosZZ23NTIgJe9lSrK0iN6ymUtm98BZwVIGc1AripUvELJPiYMozLGfTLV/mpz
AcKHJU4N6UZDKjx8/cJTplBC/cc4GibJPZ+b8CGTxPVlm8OoUAiEuz+v3+c5PuAtqrzXoPO0KN4R
jsKYDfS6aeSYPCXrUzQyCs3Th5KLFu5JT7DaIfLxgeF+06z7ixio6g55/0WdNneXrbfFBW+2WHga
KTZr7QH/joGVloHXV/xP2bPFtP0pCz/buaHwpS2ujKblhPzufMMbabH0Qi9YR8ntcHn5gRaW0qmZ
FuycRjTGMZP2ibQ98oGp7AzOFObXhLn722Xr4ruRj1vE9uwNMXQFo+NP+ed8aoK9a0n579r81fqh
N9BYO1oTSM/6Q3oi7gV7ilgfxdVQK2CgMQhJN8d5nVEWbcOOjgFDQnP5fcmU9a/TR889fLDON/IP
zwhSX4yNqRvUpUJomBx/TJnkipUsGb4DB6tE/bXajAWCVdLQisT6M+YWOYmaTFI0SKiXI1+BoInd
sM/s9JDlmmCOuVovblgBepOWrA7BIZnjBJPG99ouLrIu54AOD36SswycKrAL5HOSIWyK9gxvupDH
vCx9qt5fNLpziZ31OJ9y/H09utheZvD/4Jq3ESshvYVsDUi0ClmVMV87YxERHA0QSf9mYy4JRXDz
QexhHCCYFAwS1xtU+qOcDsBLih+BUP51LNSn0lQeg0yUpml1zt9uRLwPB0NyGn7rWsxb+F9HroIx
C0wDqfpECBFsMQ+ObbLGonrzgv/Ezt+nFD4B/b/z5d+ew74E4ytqEdnMmYyvYaggDEO4Cy9uH7Py
SOFBaEE4Hs0im6c7HHkmjwjoB2j4V9+bbgeBO9P5R72wM0avHqybW++84D5JCtxQdpbkAf0TBIlY
M8STQ7ljR2QmzHwr1SKyxAEqrVqiyrSLugV+1xShmtMK4rpMDL9JMKeINNTiu2Mf7BmryCEzSt3k
ASPpFXTev0kcE69n6N53MUsdRPETPyPHFDv18E5inwdRWSssx3mQnETe0bTbHpthgVFZmMOjVxBs
Z+tZJ/jqnfSEOTD1528lWQiymGNPyHbOgZy3R5SiJt3xWojpKPXjUmEkRFpk28DXgrgTFAafVjXa
6xXs9gOQ4GOZBZvYSUX3VWkpvjq8y4ki6ElLzkrUzQqCrdLw2KkM6IbE8LKH5gGOL/48YdVw8qzr
9LW+wCfIHQqcWyFljn+8L81A3P46NKmgR4xrQZxm6OiYORT2jQBhhJRtPgctwENN6MeB2AAp/WhS
yNSNYpu3XIwPIKM6ktuwEayPicjOK0I/VZP0td1Gp32PsRbD7KWTlV7UrxHr/17VfBTZ3UXYHs9S
aTociTCr2vPZF4EoVOyCpnEWjNz9rDYO6TI3ZpO9vyenwX+HrMN10BZVr2lNNVeODleWWEK/TD6B
BX8aUUTr4UuyzLotAleBXL8Mm5ueZz+2S+Xi0IkgEvsH1YbmS6xodZMnJEQHAridanU8gLGzo3p3
AfLditvFqok0I7My5ubLJIYKhs1AMXdyCJ/mIu/BituYgkt8NQvTJqB7/yRj7g9AOnkW1KI8cmso
AF0NKoX/94snJs57rB9rUFuNtIwonZ/N7X9vA7SYzPC4FOfPEIYf33QPVNgA37qJRaYzsLm6+BCn
HzCR3lepiZD+mqMH+uvwCI13NFMVPtqzjllpUVmr0lXc1JW/BlJ2RWoYWmtRtDoSPxqjzhaeqAwV
vJ2/FGHEZcm9SuzhXbYisDxZljZXKwwg00dxJ+Cyy78Svxs0Dyvwe0bm3IELZ2jvZxBXZxkTILZD
ylNV/NoHLkOLLlykTuGZhNyNxU0FEw+3sQMZZrOQa+Bd/3q7oXv5ltO8v63VCDBqdxfBCH+FTWkO
pU04uLJx1rH0qwua509lncwHt9nvBcNSR1iJNmoxWyzR0U3ZNVUqz9Jtgxgi7zrjKTzz7/BmU56j
4A/ExCJe1BIE8bVVDg4DnE+zniOAbxxFJPqoZcO4I+ujWMLGsmq4G4t6MCXc1QWVS4gh9EbNBQLf
X4frGocnDMPBGcs2uXM6HrFPpaBbAtg19Y7EZtQfHcBPCqLW7x39OvdA3pZFxvHAhFLU1d8hY6HV
6HTGAQk+v/ol6XAb31S65CUEO8jWM6BSsOrOCFB4QdOtTyYTElNetnNkG6RVIjFJyHvkNMqE3ffF
rveEaJ8EzXWqlx2Xiw3ZG9YZCmQUfxocKDS7v3ZgSWRbKCgn+dc6hh1Z1YoifBM7gm6JMHthTAXA
w1dXRHZfXKXBw9wNa3R3MvXsFZQpmYaMQHyI45qKc6HohVvMyXfCCc8bRxnb9Wr/3PKANqdUnO1D
VA0pc1fNeniZoWJF3dQEV6/vX8/Q+S6cp3B/DCuGQeBi80Ju6gPyM100+sZmMXcYJrZj2ZbQgWq+
pPy+D/+Tmes+t0/AaL+I8W4NDhnu8PqXpsh0xTUo6XkLn5zZRkGtE391TYP9r50KnFwrAPwPDym1
NvfYqFnBhZZhgXp82tLv2pro2Cf1Fy3yQ62ocpLz8qH9XLzpE790BQ89i42tBw9WcrXFKth771xz
SFCZAYqOB7QBf93hgE+U09vycSSPuvAwlvIPxeviqu+0w+28hkuWnCw3zBC+JeOH74LijeZYjWY1
+y7sKTuulqoQpy77DMFJwJJlBMJSBT/g4ueb5iyBtl9D3JE2TMsmnz4oB0EI8QUwCd1hJToBRllX
16KqFzhswZqqI2jxgtw/G0un7js8hqdxKTg9aYuxVzvcuUkkIbjULgwCCP2s1e4I9TJuF2aMMMtb
9mfjKxwionzzTRSfk4haRnooeIRyUnk82QMTBMaR3M4rWIOPQN7iRi9t1olnVQE9WpeABWVXpEVz
rIi/ELnsFk1ed4X8vGWxyRUSTOcNhbqujzgETnSM1V8F/QJe/RwyMY1B7Qg8vr3z2X6BTKS/mDVP
U7L3OnCFkXiU7i3qD20RD9+cpCJGINyMGX35rnHVNHoXNQOV+ZT8Yq4mFpEymQOR3kJzxX0WhSKq
BUOtn4VXTmTTHFZEjRpFkKk/L5nyOIRt3MBbA24OVQQ7SFYpMlpbVyFmvVOBtf3ACKXK5tTx28er
ntY+/GZWmeTq32BAGoC5/jxbDPWwtgUQxko5FXWgz7I+Qd1a7AvciQZpUQddLxljfwhr9qNscOcU
IM0rPmr284i25tryPITCod6l2FnAOQupWeqfd6NBj2bXu3y99h3iZAZtysm7+/YAOkzZo4BzGBQS
ifC3uH8QfrDtMfK9XnjlATqFq8zWt+cw71WHlh2cI4X7BbA4rhtIGMpgYhoDloIu5Z0K4iqq1jsw
Jbu8ZT50CB/pNkObS10seSQfSjhaPnb3GAC0hBUIBD2886ueTprLNNnQ891SCS+JMrr7NYA0Gx6M
SiiW4+tF0KrLDpgOg/tXZEOiBKy2p0UF0lSciCG9s4WvxSiS6ICeBhmlxwepKB6VY5CYqSC+09Nx
ZotklUmNbE7ljFkDVItLASaaHTjrKEOsgq3sl3OfJnp7C4TOP/CFK3eRiOPbWqnrLOxNhzoIJNoJ
le98nLw9IkWtfv9PpwsC3Zr4dcfmDV59a8aMzZ1zyz+NrUuCfZ69x5ma7jfFaTTBPOCMGmlhYhsu
ioDS8w4NI1VEKAB4A9ieEGyEVtVVVVXMZHKPcn1J/q/17F7qwbLktGdowFkxVWXhKfnW+b0mXblp
FbS17U9n7OIdgwnO6G78tvqRJtaQSS2mlhti+qPtikH4n+UrlvFs1a+lfKfn4/4Ucn5A7mcWkNsn
ief4Kj9MenrxHqdoiOeeoGWbafL7KwGAQMxv6jfUEnMKa0CX4riRkRMh9Ll4UVeSQvPunQ/TsVag
oIYkkV7wugtnUhnhU/w3dvhuEhwNO4NiJB+MehEQCJ2G+9L1DAfShnZngFMjTH2PlgJEdrITVRs9
UrXf4LaP5etdNo45l2xDws44mJMh5SxovwaMyx0EBgpt6CtKtv7kq1mjNkxywTnodEuF/4Dss54u
9vE5YYNjoTdEvs0zej9NlHC8eXMdnnZQmi/Kg5cBKckZ7cAsw9o2xF6rjfsKuObqnIHN5B4RO4Io
LsdYTnkgKbLz77b7PrikbFxdJmziD/AYqp/F8lDXfw0PseM1anQOY8POeRXO8owaGSkYsnMqeWRI
yYnUN2uARhGj7ILeqqUZs7EIhl9PN3dEUtxjcxzYWQvkWrFjaxJfYK+12RImJ1Hcpt35o8f1pqIH
nWBYHO1+JzFxg9ZsHyqZSAYg3JE3jbNvnGw4zsbQZsuSZvm+RGv+95Ldl8NoCKm0PnWGQGDWhpc2
bRuusJ1QIEP4agEbqwLPoBYyb5/N01RsP8WdIFmbMpdRQ2M6GqEXQgxVxuTmrsMNeusmuvlpuunj
uI4pRo8B6RboiUKDsqHWQnzMbKRQv+njm80XwoKTgSTMM0AFrIs9It3RAw0E/YDyym6vWAMjWX3N
HZoSLg//GU5eHPj6d1dGxr9sSekX+O5LY4iKlxlM1J5miUhmnDaxjlrAjyJ/SHUZbHm7iE40ZS19
qX3gY9w9jW2orVTetMi69GE3UAE+bh7ju50BvZ5gnfnmbjrch7hXuDniI35MvGlr1UigIXcTV6pn
lZUg8KTM/qeUULYwbqLbtOyLY4VluhOg0CYX6tdbrSREXbGNMtJL41vA3rlAxw1ZKghIc+H2z713
B4O8FmE774TlNflLWForOpxyy2U411R+6qFHbaMxn07Vv+NsYZmyIgixftph2Ab4O0r4fyvGuwQW
b/vyiOY7Wlm6toWaMSRzrp6u5JPeENpq586yD7QT7Uury2Bk14P1H9GNlSq46LMCzqs57YGN4dBO
ki6ht/j8UUeGaf7pF3HNv343Nlt983A6bATM10yxLqHGnSiIR3c9UOGU/ogtOVdQ1OsT66/74dwf
e0orh0fL32N+9SwgXfQne7hHQBsagzbKA/bis6iIrVeWF9Lel7eWGeHz/RjvgvlxOpD1NyllxTYy
1DdLcV4iGueiGFgJ3oL7gbfTEONHjxnrrEUAYEIf3QNWKV1LKrWP3YsOGdz1WtBux6pe9Nq8sjHO
yzdoc/f74ShcCsANci5Teweq9vX0pBMhHyO0Urdl39YlTXlkfFApU1cuWYvmLGlgiD+aujiWAoSw
PnEYhHN+Ly9H1wSEY72z8vkHq4mtu8V1liC2xORI+jRNulzjzhjF9otSiYzmigLVuaUfAgMOkyIG
ad5BUBkUepCkChPMzZM3twkMDU/Gmu6Iq1Koczd0iIhhkN0Wdvl8sh670CN/uRkhJT9v6nDRnFGA
4dYuogJRRTBCfjRiWahtfI/jt8om5iS86ME5/oyuJqcJeRNUXWc7YPdQ3EWlpJg2KJI6xipYluKU
POAqokJi/PENQyzV33rg2vJeh1IZQXJM4IRHc5k6hbLuMBF/H363eJjiqe9bDw+RK/aEkrWg6wg4
6u5lzHjW0L2jMv824cJ7F3UzuC5qu3d34jHWAkfFt0Jo914b3T84UE/2K7zY1cNaO28UgoEJ4Q3l
7c56fdr0Y0UVQ0ZcPPDSCapvzr506uugKnT6Vf9AfgWAcTo9LbtjF91tfrHADec6b9O6Q8lodN/K
liWQAmqtajbjLoyiT6hX3adnfMGpRJ6VCjoiyIw12BPu2yTbxzfVFicTJyoOuNrUgzqBvqNpmMzu
0kzgsv/xUnotsoBRC2tkS0nuNbPHBfV3FiSoT3SoTozf/9+QB0H2JKhAEBO2H0zFayGEZw4ZSCSB
mfx/lgvc+duKxMERZS4cZf5yHmDOkmeU+ZF5WgqDvwRLkalCPfjDOkr2l8Jhtl/+spBUBNfjM+Mr
t221HAuzem0dLNktHVXepskIkshbh7c3XGfN0midsCW7NotEknFI4M3ZFRHxHB/VMsyseK9VZ7k0
93ka0JzYuymKC/XEtl7YMqLtYOcnZclUC4z3kZbdIOQxRy1qiSPNQKyDnUx6X3wJwZx50Rvtgvmi
9ifCRa4r2CW8OIe3DhsB0F/AFVXYu0wpNTxVucNyg4WXStBrrQH3jKgjXfcFVZCPFPcfZXMf+e1p
WZl+aU3wbqIHhD46fV/BGrxNEQHWbeEnEdQLHtRmoCgCFqurqw0oJ0X3/xRdtrkpREMZjCe9T7JS
fcAt+hJhRZKGYyJfs13SpPcrNiFBvIigatDGDlVvhDCFKGlGfEQdCoA3djsf7oOJ/Vz8xkz0V+lq
N4zGeU2KI5d/FiXjg0GFtyfTKAnG4UYYMjmWJUUJmbmQoXR3+0DZxw6IM+FfnfvApuLqpavBJdN9
7Ku/mM5cuURXcQPDExVa/4VkI64W1Zu9XV2NmIVzXye118C1qFokkAz1a7gg4RhA1Iuc1tYqPso4
HK3lgGa4KaMS4t4KFSrv5G/A245IU9p6FyMWpejS2QE/sprHn3zCUKVZEk+UAqiBJRXGnv7R9hI+
4wdChnifd7RsLMoR0xDqIBVLVd3AICghTg6RbFTyQ0D4Fia6pvi+hz7dK+/dXzNAi86yuwqpDGUI
kLOerYsv2m2W94aSn7X9d49ox0UtxsBuQYohjruL7kKCBPS22O0tS++xeNIBUNvp7ElMN+HG59O4
Fejdolw7YBbKPfD/RZXGoqo67DpHyoNUUuTtUYtxER8tzYCblZ1EQ036esPjr36wSgE0LdOUendf
c6e1Ay2WZwv6y4ZDf8eIfxLQ0aX5K9zdt+FqjFeoeFphu/uIL4HweYpvHzckl9V2uNLJwCsO9l9K
iS+T4Ya1QjxzUrDU4OQJHA8OmDOZcWZtUohAi3w/we6VLUGzCDroOHy/EjHSdEi0nAVLIjUkHDep
DVgyAJ9FvGA2NPzWE+/jTXQ1A735lw/scthifOsKivtASlrp0JplgG9zYl6JBOZS1NKBwLcgXccd
9/dJJQsg2QBoXPlX3tDT5T/mTzlyCqmVplEaUcVxND+W0ew4XjMkxdr8vIXMcNaWjzMLxTtdXX6i
4sR0iGx4ZkLRCNUGN5Q4UZYG9eaXq8fsZDzhoo1y1GKJLbrO8Q0O3jQH5vzd+rKqjOiY/V0ihc8z
2knTuIxScQD3bxKrPtkCxl6BfuxUvKK3VzKlCa6Ss/Zx9Kl9yb2ddDQxKNiRoAhYZJnXY/Puogrn
r1ronML4iVLonlT9A7sEQJwkJBOktnrvAM+GahOVoY1zt4/4p2heqEQcIZGP5vsEUxKcasernU7/
/1e1KWd0av5w8s5RrbnVMzK+s0ppdNub2u2GQDKxm0MEzJ+vHVMQ9qEzxcMkav5T/aMotZ7oPHPj
Jol5rjyuEYBckaSCENqx+9MlGWU1aw9SGKui2uZsUonAwfQJGuQAT4NxmD7wZYUyViSbw01EzAlf
W5kEJJb+OftL0YAXiMppzsLuzLVf3f83hLqdMlUMrAoyDdu6y+YVvBfCOT7rCqxi3V5XF22HcCY8
RiiMOhQyUl2eMosftLyyH9SH3s3asHF7cRxmu6rsYb954GsShejtTfr87o9LlnysC9SsVmG7jl1k
UmyDIGnca/INbLYXmjHaOhFhcsKMm2W3qyKjob+LZ1xUI9RRAewntYXNN8qqh8dLXQces38J28P+
f2NmrPpOgEgMpm8lgUbOxPQYSo9zBaFYqbiyrk6qgXN61Tan5upBX57EYduCHTtz0XWykYVhK5Rx
BNOW/PuBCtjLd7NONljOAr11LZmE6jXB2oHK25xNRAhkL42kiX3ljY2FCm1/gxpe5D847wRc/U4q
VAhV16HkAo6wks4+YYlQuVO3FuAytvDUlFpfCIm63orcJQCgDAwMdhhLNecUDU908LI8BoWVWGls
8pSGKU7vzrGT4lKO5mJM1MPNMCZubd+4mgvD3vbD1vUDx5xZMKEO1rXz1IzFmWQVOUR3vlO4ZOz/
fOaSE1bj/XFaNs5akGswFih7YaJqzAyQlPkmmIR9ekvROmXe5ZiOKhtRjmuvKhC2YuAudGyBrJN/
B1SYg5DxiwltXKkxROx3CZJgIMvj/JjQ+vDzm4uGlYwxnEOVAIoOQJKLXXP6xVE0M5fsfk6iHQCa
7NIP+aVmNe7rO8ONQCc1EbxQQqNjp9C/87U577o8gMxYvZLwXm5QsjzC7OOMW7w34Xs7E1Y5KmHq
tQH2g9ojptsd+OYBa81H148vqa/wf44EHKStEj7QmwiFg1KlzKkpWLoPwLzKqnk4ArPpHRThJgDT
DYMKuspVdLnIrcMrA7dUTCNa71UfvoflTdJmsvGzHoPZh4tOwM4X6llxDFmFuNrvgoAd5k2gtI+1
hdENPLXxAmaS9hONY9216Kzlt0sjv5AwnPW5+3f4DspPjinAxsarDL7U54OgFqjq5s7q2Usr//vS
mnm0TNzpSbIrP57SXXFeF5MnXKH3LBDFDt560zmnpKHcEbZtZoL5mJ1ipjhAGnJSR/wdNWJiK2BG
zAc6UPlKxtdyQCzbWbRbbmXE0QxO7q9jjtBpEAIMa4LQCg8GQ5ucWCS03WZvVHcy97WViRtnntCY
x5DMAaXxufZ3pHHaNeZmzW9ZiMxCs0Cwe0pEwPwt9mRAMG1aEKrIWM+i/1Xpalcp2Eb+nKuBZX14
K4CmqNKlnP3di2wnOCwQTvJ01STIFSceumGwd3QiT5dierkmgH7ykGykSXprec2f7n6WUIWmkLY9
FPzY8CvCJPn9WK/6fjEW+G3ngwPsa6jY81XdvSFgqyVB9Xqv05JtBJ6GChvG9b3GzIGseMvfFW1d
rGmeGu84cQEDlyGtEuwKME9pBbCWnprmXso6D5ICaWRSV8Cqkrz+T9LcwmY7yEw4ur0Iia65Ftky
lhMDiMPh417fwR5EePvriFMOMhWPUaHdrYJS1mS3Ndc/POhxXOJFtwaqoV+TuWD9O9M8G1WGVOya
vlfAcZJUTw4Si9c0vi+ICDrXYvO+edpPwxz4Mpw83yGloTPbG0nymuIzy6hcdQdJtFpZ2tZ2Q/qk
XxB0Mw+CyHSjYWAU4D+YSwMgQM1RYC7Jbd2KR4pM2ozVxvPF/rtkw8Pp87Fp7O/2YPTjBmulNWtD
Szk1CFOifrfhbgMYPQFb0KJqRNvcZ+L5nPMAfReB9HdlA8x7ZW2c4MjDa+6EGwX7ot0lc+kCujWM
KNJySvwbJNlHqpiNsxMTT2VjLJTO1HYV6kI2jKosFNlrCm4g8k8h4slwVCENlqZjCEakxieSVoLI
ZNBKjyO5OMfACcKVlSgqh0RRI2F2r/bkKuehMeTEpMUrneKJ6NmZUjyiuBI7WIn0RJ7OKtUTEMWA
wy9PjzmnzvFGDXk4+PuTmHKJ+u+AIyhY9xUcunm9jKBMX+x13BHe//U0v9Wix0ajkfoB64Qkhg4s
utcZqJdpYqtj7p0vsE27Q/VQrKcQXyOj09J7TpKYK8QsIYOuxg05qa9SXOXEo2bSaJfL92YsmKin
LJngotO4wiO1O+0H49u+0xXzmjoHAJ3npWgFxtvq+XCSDZwRpnCxBrY+kG8S+pL3+vQS1h3AQds1
ZBPlIUsKkTci3VwkzvKDpuqDD1ywwd/voEWRo/WsCObDYFQBdbufHThYNjx+g2dFmnHyFQ0Sgtf5
Y3esheAbI3FUYtaM2BMmscX9WGAySCUXw8rh/g8dR6lCQC05y98vgZ0ynuT7q4CgIo6YtekMMWvV
NYAWy+0RsWH7qfETZ11Du8bfZ+MkqIrsbGpZfvUuy9PQ5dMJlrn4kb3y2+gFj3yyDrWC6wxSEhmZ
nL/olzFLy3XwSQjlYuxOnMg5awY2gF4z6rNbRjJ/DAnKBPnwlBsrEZ+omvuaJSWIgengqpqnMvNd
z9gHe9vN0CYqHTdzvtH3NlPgejyDdYBHYK8vTteyEiyJwgb+vE1LgLD/Grp5dDzVvtenzfnJcZnG
OLvGq4WMkae7McwpPEavJcCj7BQW/TxKc+/0nsR7EbtGMGtCu8OZMmshXmQwuAm1Pb6d5AIJ97uY
WTZZz/S2+Hf/mst/QXJJOTHSCNZHDtP4caymkIoL6k6ju1V50jZz0s7FXmOhLk8533olu4wKDUZE
LM7mf+pSJWRSVmbvK6WWrECgE5NK8NVr8o7hKvqwF6cCdrdSpGdctDPy65ByTNupEs5S47gP4Jak
FkJlBCBwhpJqvYodGBTT3c14+B9M2ZXXAwf+Osj5Y1sc/el1fK3c+W65H4YJGhzI45K/TLGTuKtV
7qf6oH4VkxJo4PXh6245cRlzdmXiSGffA70I30B8cdumu17VnIM457gP+sUNKxsndfgJAVw5SU5Y
kn3sju/OFBHKvX7FA7oXUIMoNeIoloCrSB8eaRdTiWb23rWSf77RHtdx3y6TARn/wIxVzZVOnfPl
G70rw0WlGm8OaXmnIIHKSl6nq3jhhf3GpKtKrHJwJS6eetohcEsUwKIJT5q82SGwZHNAhbXaLnQS
mIyvyklpIRWgELBeosr7vLAY8vFmUyaNQc61Bz46cC5pw+fedkzLKm6abYPT3zjCSqy4kyDrm5dX
cozX/Fqsh3yIAQrpNa9a7T4YlswTqm6XNhCu8wdyAUoh2Zb/nQ8mu1AUYwYOCgF99itdm27rP9lK
lbgWdZeN8GmykK70i0ye3o/CiEw2xxERN2fnkeBGBGy1ua5/PloLAoIhfBAliYEWRja7mZz2cqXV
2mHjQyqnzTv/GF1+s9ZEQ5hpTXqbDvhBLvMKVWmD3vo/hxefZyjgmeTHTC3LQw2asdmedskyV454
cOWsKjJQWU2PT7L3WcQYS03DaBvjxwfPKbgNUo3UqmySZ5sCnCmB5l056Sowrh5yMZwZZr/DeyQL
DCzWBN6PR/Hwm/XeVYpG86gKJtKWVrdsCZZZpjYdV/Sc9UW8DIHDG9xQw7YJv0sWvVMfVHVUaTs1
8r6DaTfRcI8qsOGGgtMxR02XAlmoba5JolmK6kjnqSqAlCnfSz6kV9cTKYGlYauL6pduKryGpRUV
7AfY1y/JSpJ5+q8P1XjB73ADtWl0C5pB/EindqnWGAAaF45ezyiBw88m+Uh+8TBeBX6k+5/44xQb
pCVdz/4Dy4NZflbPIEZ8rqUZ9YGMGKUrF04Sx491SNyd+GW+F/nghC7DgZkDpr/qqRxzpQTwqM5O
UB0J2je2mbgIV1OKWi0dfNDIoIIeHT1/rowiwu3mkQjgMLqaoY/aO8ORHoeWEpCln1NC2iAMoo3P
LeQOQZ9S5vcvgjSIpcN9WH72u8p4MSZtzKu2zK5FgMUaBBQMCcgEkpITZqB9UHrP3iZnR+3pEhZ3
cD1iLhCP64sDVR5+qri3cTiDIoPkr7HLIcZ2Fv9n+LnKvcyoLWPl5KQTICP0/P/Ad1XhMOeu1G4j
rDWh1MVFY9WzXc0Qq/axX7F3pcirQqN+voBVTIjR7hHPEWUavzllHemvbiVk0rdpwSCrs0FB2kGK
9GyB15rsmn4cuVX4TzVyWB1AJrvB/Wv2WSPTAUhE1PydrII9XXl1ZjNIYqTuRaTmTPg3CdaDv9cE
Fuh3cs8gRMdKTLX8TSiBvdMl8OwOr9ARWdeFLFvyVjUnuL9xBao6jmKFrMGGyDy8BhNj0gikfjRA
piG5JO/6JT72SFbD9Ij3ql0Msrgzkqs+MU11CMVpfpdVapv17jd1vYQUXsG7ahyVJZeKsai89YBQ
tEqVte0slBqOyocyxeR8oPu+zLXvilOeCXA3/MphJfMpAdf8ToPwbVwASpnr5U6D8deCIHblFAvo
iwbOHGCUz4209rUT+xEDRnDlhBJvxhKDgFUpS3xshjMv7ZcHahL3Qy72Wxtpf5na5lB5h3IkdGBS
uMyywTZrbA7jOOwa/6B9GOD9CGQRkR4wgIh+/XyA6PdD1xJTuSTheTAsf2D96ca0/yI9jvTDasRs
OHwT5NHvzqMBqCmeP18DMgWSNSdRC+ZLxgaOSgSHE94/pNil1PIFOM9rMikre5UiDSTBadUKcKOe
Bg2Pfg0yTkel2j8YN/f5kPP5mFancSN7vVHi1FFqmxd7Hynsh4cQhean+ZSi9rrTbYhAqeFTpZ5L
PX59ex96bbTjqSC1desaut+sdQPxWnyTImX8uGCFGZPvsVcS9DZrCCphLBfGjQ6vzxVBUbRl/xSR
J5QqlUjMeavDb7pRavtu/RJ/SvNBiY7FMTr423Hwc88YUVCfc7jFEJFWXBsxAjwTUcTIKBXJm0jW
08pI16WdUOq3v5AjmfyWbTRiaZRxt+sPiGokRxDDUsXS2XApoOHN/ikn5YQJuBZ7cG7yknxqHfym
jyR7D9l9l0mEV0Ua+9vDVrmpcK3TASHyPiNn8rxK798xAT07mPYn0TRYxRTarnrSLQ5wjwDvlCzY
qDYiaiN/51C/Q9I1CwQyElI1KeApkt2wD70rQRL4819WBDVZkmCPqUTuULVnvkj0tUx3P+/L7qCO
4GdDXEvQjudxJemIlAYRKSje2GLaDkuv0c79pZHdpnBi0/VKeA1oeeYjS395S+tlHTeHbbujmnxL
vC3uPI0SiHftLHO0ASeWIFfBe3NRsz7VfuLoBXEgmRMtUPBeP/eXb5cua8QA/jJ+2yXYp0CB9HN2
GL+m4JADqaqB9DYOz5MjOwbCHhJx+MMY2LcXgprDhQTgfvaclWEgqatt37kFWy2VHTjpYvVgEEPQ
apk+DqZw24B5Cg4iwxMG5HCo5isZXaOn/xta6F3NciZY9yGrWNjUvHPJRrdHtaYoRjmHnhOs9jz3
nbxrCZd7FoarZNCTLFuT05b/W0JzcHeN0a0POO2SZ6jHCL5bfz84Nvkz7WuOCMj+VMKHZAzhOnh4
vqeBRIxhsOCCIV27mRjj5lPtnV0dvuPsAkc6xh0i+tqbWTc9Z5ikGjq7KKHchUVHaMLCYuocdh7N
ULNEwTk0KpGR1nPkKxvB7M7/F5plEdlBbo84w+2icTMfVGhC+MRk/4fYITD7/vw/2TtvSUQL+UHo
eG4fQ/nbSGm8be7nYPnE7+6zq3Qemkbf8/vtixhHBgItktwwovWdLUKelJFsKxxWgbqTamD+7mX7
H/bfj+za/KXZ6bQhqMZr/f6x/206ZIR2LLwx/avVKfPscvnx158r6XSyen4sH+CQjfAffpo/kJNa
H+tuFxjI6WEioJ1fEG5pjBCljsd0Ahk1Wj45nI9r/dkChXs1VSVoZQk1j3uv3xCbTMl1EFY2H6h4
of9cYwbYgJg5PJmkXx/UTzRa0mLtbs2fsvmP/vARf88hxxWpMu9BA7SAUyrCd2oXND0iI0FOL8R1
BGq5p8ogCfGeP2AQyoMRAVbjBA6oI9iZq4R82mpNMX6yCF3jaUEnufFINpxz98Bv+IJcAp1ByMFD
ySU01l9OgPybusp5XQJag+ZHgKdbRQX28D4LquqcQ8ycFHXf5zzDtttTnx0D67dFkFS6UuRnSOef
V1KCVarz+FRlCezMm3fEpOvuZWDOUdaMHl26fi47tP7KP+nPENTVVKyxrqDalDBjItGQA/3f2MIs
zuqDkhYeuvnOZPwFK7ewnYTkt8C3GfZr4aK4iCnJ8IpmmFELdrLCAIwuTMlv+kEWor765JeEvP4v
IdSco+fifw/PNGx/DlrJ9U5aKhlYDT/1XBFCgHR2mzOhCszOSN6pmrDMQCfbYc5tDKDooM6r81xk
dYrq3HfkfQljX+e499gGs7FE+7oZZH9WKXYYeH3+vsUG8CTrGdnPxgtqWf72NXMGTXKDGII0BUFZ
gDjlCC7h6lIZ8FffwdSicnjWQuOVtxOINzJ1RVY8AGrFYNNFmmRDZavhVTRV5LIodNdf1rutRXh8
AOYgd//I33oBcRtShHI2gLCh3OuCWVHb+riHtLOz5fQ5nIFuzhP6Zdg4Zhw+zKiWcRzBqCJ21o5s
p3RJQjQ0obMwjgirQWN4R99LhY8aBjJJ/rvkd8FIgM0iUIPr97UMBcdMUGn1mDzvxEUIsWEepskw
ebvU0+xpXEeVmnNBmQ3wxO7AOv9Bt3gwagn1AUlgic9QT40fxb2Lu2c6jr6lg3FeSZuKJg/R/b8y
0qkVP/0SLgcNUV+gU59eW3IEw85t3fZyJ2wp5dpWZNYvJMbtRxpQTKHKuGT8Ozb4Q4Xup5bRXKPD
kbOHaxGSC+unJEuNdvCLvINtKbVDcZcqgx2KuhA5Is6FKyVtZNmWX47KN9YTEom1r6CDW19Yo/cK
jBX66X2l6e4luWuQQCF72Fo4C693c1OKb925e9FZW56S4l913yI+Wnnh1bkFVJt57uIUHZa8G1oD
45c55oG9U5lwwcB8lzak+eFiO+DHi4w8aZ2LkiaUrlbvLZLu+EEEEFNJ6F0j18b0/qW4FgWycBeA
S+ttHzlTYhOY+LGW8jIFrg5FzERwmr4lcwM15lDkWHw7iHY+Pr4HwTuZfe4WHmA3aZIhG+aYUilH
sWmVpe7Vmjbn9yCrwkzxK7qVaZCvNafCDvbqIdD5v4MwjFHSgdxSmUzRLQMLtgkuQWorZejaUut/
AUu67mK1NPcNvyAQ1cJiP11yije6OvKvX2D1DbiIyfGVdSOquJH0o2z9jXHeKb730OP3yk+M4pJL
3fWJepszBAuBDfyeWhYBkgn96YX0IDmLLfgUfHKFt/LwgFDAnwIesaUY1pVyYeIiCBY3fnwW8AOX
l1c4Z2UVChcKGvVqzD+zX9qGSbjZcyugMpT0dSoEG7ZCSl2uDZKIjQzM3cPdJQuI0KpppJyTLdtj
jblM7AkVMYHjMkWMl+rvdd/E63tKozDCbwL0NpGiwsgtcU8eEtczOSiuhU0gel+TkLOxZsHJqeE/
f/mAJbKvCG05XB/tt73/H1Yutmk0rHa0j8qG40XDCfDYCcKn0jizaFoV/qcHtsn3z6H9yMpKbYoY
YcRVH6YPn/KayT4TgC5fKSISxqSsf5oC/sQwAJc5UuV6v0SiKyEMCVTvb6ClbyXhJslJy6cRAfJs
45j+PZFt99RgxnoiXTxFdPToL5nGPgPaElJRAiz+6weX58IYzY7euSV2gIy86hv9iihOsBJ+VWAK
DJtHqSfgxIRN65zKFaa+7aO3cfrn01LQzBRhSNAvzAZVvc785MGhYCQb9eI6BcxMFHEoh86HmmoU
I5CFsqu7SJvLDjwcRyKI2QXOLmKPKbbQayoQseWfySIgMUl8XapEYs3Z0+H9EW+/1uRjtsec92nu
Wp8NHBi1EXhi/Hjvfbj1WozYexaU5Eh55TJV/Ne+8ljqtnDOXi2kAyMPaMSwJXvsL0s2h52fq61v
Ycn8+NWcf0D5YSDwNpQxqMfwepE2bYYFGy3rdvhp9YJzHOf7GdBcU9RSlTvZ9KBr6JZRaWQg/csk
7USNGQVMnI4iQQo4N0vnRDfMgpJB07W5skusj9jyjEQpqctBzqZpVMHcIVoGQ2zeZvH9SF6t5BCc
8FXiK92g3gYd819EBbM+8gi43cBEiBGhMJr6Yyo2Pq5bW6BAXU0g/GMBhjRZEpd0vMx9npo0mzBl
rBjzjpNSs+3/4hyZ9hTNpIdzNm+GMakrcdey5nmBHaGCST8jAW7pn/DO0FuuCwFziLGGKvEp0AVI
BYlKssFrW9fQQb3VcpdEzJN/2Bww+fHbrqC8/O2wn+3P2/xUyhTtYZRSvmBQ49vbbl58cO+ZVLOE
vY3NsoaRSIh4IG2T8DMj/rAAuf2HDFfeoGe7VR1aLMfYiNNYBFkCdFn8W3R7RVRsvW15upciAcmW
cgFvDX5ky51lJYJh2Qy0TKa46GTTL9fxD6C8nYDEwX/tJWIR5UKsKIfk3j8M6wALEx2fZadKErjY
/n76Oj584M2pmvlImMAPDFAH8I7wLP8+1jvUTSFzkzRyn7vyUD5v9Lov6pOKMFXgPtTWeu2HTJWR
57ICsmbUwY8cYhKFXWMjzPLJ+TY8N1vgaz03u7HobhdWDncqOBHKY6ECsWkbDBfZgL+8dgjFwttg
CG38EKOI2jqUa3DzaYnS+H3s7y+a0QsxWq0U+Lu+S/5BQkq/AcHaQmosPwgsfnc9P9UN666HRD3l
p9t+X5Jp2JZvmBlPCPzIDbM2k9CiMsJwkGCxR4HSy/qRu1GIK/ha/ufsGjUJhrbTwRT0zxRMcYb2
c/wlqM03cv/AmjHxVHbCTI+0Tjn57wztOBcWOjMfZTr3Oja+GGX68M6sxm1MZY5xVDixWDPgr5pR
iMXv8r6BVoHIqVUOGd6vHCVSUvbaa2vCdF+M493h+zhIKg+bd5X9MDRHePD1w7ldWCIZ9e6kqgx7
Km3vnlkF83g21rjjvNk6Qujr0gcUvEOZpDJFpK8jti29RWJ3eiMSpV3laYZpBjq0V3fr2yINDoSV
8kKFV+vIN0WROKZtT4vDtYIS7o5r7+Oo/ZbkwzfBtM0ug7xC9zmYCjbGC8e2BTpzmgxAYOdOOwVD
C/0nPbdPAAj0oLdkOqi8IpiZNhgXKV+UPfWJ5YYIRrgOVKFOk9wk6euWZXWLy/nuV0XSWhN0PUIS
KDe2PiNhH2Qa84orCcgW+HyB1F8A/NP9DcxNajOSeLa2RTziwPD66r79H0Q9TcGGFHn8i32JtAn1
sdcYql8eND0GdalKQSHQJeGAXG8WIGkBY94A3i2I2owyur1thRiS8RYmA1CAP4vZyRWzFzDghUru
9KguvglJTgvtTzdF+2SmyFqmyCeAJFLaLdJhFOe5QK03/JY6Blro1S2L8SXfR+aSgGa8TsgX60Xs
7+anygznuxXHs2rjX8TplcBhPSKNOv3+dmx2rDWpPmtWPvC9UFMQrye4NT1BCx/JORjBfhrlPpPh
xEFbK7zaimVFBcALskVCeuPXVvwN9t1qPyKYJLZb8JobsTtSn7SFXlbT11fT5jjjzXXr48wE3D7p
3n2/JzXKEbabrEJ2PHxzvZcaljmhmnOUhdo2RzXZolFW79vqSzscBH1Z8fQSGMDUzJYIzsZ7OQXJ
e+k0iMY3Lo5tNEi7XDPsjwviQ6MrydRkUj1Aax6DaFA0uY+nFt5XzKxkgvs4rS41r8fVd8A3Jz4r
my0mnl5wDdnPEZh8/tA2EF0e/roffeSYNhrwbyvYcNWIHanKU0icHgmLfjfYsWnjiTdPzvrkYEp8
xZ4G2B5Ny/DD/npD1QXXap5UvdDR+2Ell2ue8Yxc/xXufzXG1W3UzGlEbxx1b8KBYIioWBuJtLNg
HDkziALMBKZ3TDd176tlLytDv3Bf56+V1FkD/kCAxvOx9PDuVTNkclUxic7AriJ8Hc90vDBtZ64U
SdBsEGBQFZ91pfr3di1zQ3k3Ze30wTBfsJuskdZAW+GE7KAlpkRANsdG+nDBQS6d2dUgITWf1Qcr
JByo8A2q6STYbovQtB8q/1O2yyoGpKgg13s6a7pYOWvdBYvPWNfD+esuSfxLRB3KKhr3kuYWtfKy
XCNk6fD92pLUZ9mJrG+6Bt5/hKJnI8yuhD7VYydosVlMzbFh1c1R0WFhaWwperIDmMklqQ45df7b
bQIJEnnl9+bX1FZ/LzOM45hakcdNpYEsgLVz+3AdQfnFWRTfYy5AUfZ07WAV+uAgTY/utNxq/iQl
nnd44xO+evYZX3jhlwASuc6qG2x9E73ljvym09kwm5oiMNeLQzcAlfJJ/sb0wQpZtCtkA/cMGAe5
2u6AmxOMhfkdPfBNA57vQMxuVFBXY0l4AJOT6cp7KhxyGkgGyXFCJR0ha5izppkA3G3X9PeltqNw
eS/3UYt9e7RWvP1yI9F9DWe6W+agEfPfEvqGS9mKgDkVmQQQOMisv548XuTPfpASJOYjxkG0M63P
+3bM43t0D3imvt3HnsuLaRJfG2c0h6lE36HeWUg0+7MLy2JCsJSVtMQksqmrr7mucWXHlGeb06dW
i9JBTXA93kbsC+VJgvbFhpwMu/NSwziLNn5Fl3b25R5aHCLlkb7svQVOygj1ewlUKMNC1zkRwNjb
c58ayV5j9Jw454wnBoLyWlbWfvVYU69X9Vxl3Ti79aCygpYndI6KdEDiQtd7tSyHdX6GEOpv+j8X
ehjIz8mdHwtd3eKVql1+qrOKpj1XoldHe119fLML0nq1REXzqM8ZwAPNWB05KyQD2ZtB7JI40ru/
fR/PNs+aAAN3F/OixKDD6NGS8S0vpUDD22llwa7VRxQL6JgC/PenqnlbEUQpAJATpPZl5dXkGWBG
2mUyy7rA8xIn0E+THSzLBvMA/WgM41LyC1xRojro+t6PAFNzbrL7nb6N7FIphh4As65hT9q814gF
UDPozPi1IC7R0epYnA0ZjBkZJIzlq5KQ7ePn+mTdgBPC9K192FsSeaHv4rgGwXo/bsj4ap2JZwDs
9E9v9dAsPCBUwx5dBTieSVbz0dHJ2KifguinHq407mH3C3DA6ThuQ43/N/KXe7CtbqHwcmjv4VtJ
ZVi6qf2My4vg//bf9sryNmXzSj0RacERZ6QeR/1iz+X0FS8NKZ9oFhHrP8MXIHwsktbWHaP7pR39
4kHh1P+IIqYcGw3PpGBusX1w+qdLBEjY+O1Jvp6fX3QedeVEDC+4jufqKajzHmoZpW+9R7ML2Pqz
CTb/zPQYz/QMDnWNh6pBHIZ+wBk/nl6P8iwqqg6i6pbAHA7Nuegjjwf/9+ZPmvRp2/yY16oyNiz7
t4QsvI3IiV4qyy4ahmkgBF/KdiiWRmvD5wLxagdkEo3Nldo50LrpTjjddUHUxjjtglfV6JRJ3jWO
SQJED7DVOU6sLU29qXDthfIu1IUXkwqpappAaOu57mAE6hN0nfXoV2VELRzx01vaxn4+te3cOecn
Q4Kn8tSC54piwGYQKdCQ9/ySagAVYx1EPO/g5OY/QOlvKRDVPnzGpa8cVCqDxQonxrzfLAor0UzQ
CB7zN2Q2BzFVSXAPuZfm1fkI7KKt8/K3B5BAuUwnqBshx3nDHF33nOUTrcqsn5pBQggCTZyK+B66
RghYGHphsuA7Fx8Ic6Hy0qFb0Z7JpX/8+MU0hVlaJZYuOquvTu2SXAghaSxAJpTRKjUFa8XbV6zZ
SZx9bz2LSjKFjxU0TLdw+Khcw9d+EruMHlbS4HS6QYNVjrotOeRvKFoiOG+viT/URGPcU0Gkv8QZ
VizzT8HA0zmawK9HZc6IN8yCvPN17IbgVCp2fnousmzOaTr0O0HQdIvnIMt7wWa8pySbS4tsHpda
nbLIVjHzGnxgIHGXvZU6ehOudkMwYbAzth3uT0D+XM9UfLwhoX54oXp5Hgx+0Vg9Ri1Mrvk+A8Lk
NB0ks96TFB0zrSqwXaNORqk0+zy7HhsVOIEWzBLj1KQKmuuvp/eG7rWkTnsRl8HV2Jd6fzmRAji1
wjeGNlfonIJWMBMYbvsxSqYPAQ/KHJitdF7XZUD8VN4JjgFjLT801Cf6Re+qPAhZLfcXjmIBybs2
WHZDcMAR9rRiR0pOa7dRlbCDuCzZlNMT4z6/73FlrPmaJdpVljBXjih5ZQ81SmxFEZNcNGWykeHL
dvLHbtx4jrxSbXfaq9ZFxhBN6HzXZkg+mlrQ7yb+pulb/6dUJ5hN63dZWkHpIfN1cAL5OU4ihh+J
p2pkVXoqPS/nimSk50zv37eOhfCP9nYyQLMH1OnqHXP7tMuE71n/QLP8yqbzxRe6uIipLNMkv+fK
GyqlppC8D30Bl/Pw3f4XTji/gWWE9uv0csRfKyG7oJCZK37bcPoOPuTU6h1K6tWIEDsuym7RWF6C
pi0VGIOHcAztxQHd1TfI3bbPVuAASPWcQhvlwizQbvUdUou3RThbOurYrgf/C17VvIpCIhaz9WuR
9dM6EOd1KFPrmA+7/7jrKr0aKCuYzFT9ES159/O5nbgc4rsZZDhcK3XZN/kIrPex2n2lHQgAughh
paK+c8cIGxYjLbT8y3jnJ1Z8UEM+hv9/LlFDzrlvYD4t5dEMTgllyuR2uqCttNZ1BVoI3/KJwwEi
3mrlRUAfGODU7FvrWGZFHDwkCVrqNuxU0yWXlXAsvntIV+MHc9RgVK4eqtYraM2Z5WfW/BOixmyp
WUyNUaKx2RkT188LOQncq6vCQXQJMSWw4tvT4sodL03D34CtYKnGTQsxuy/JEOsktsmP45vGoSRG
DG8vsZF2gWhh4fMpq8IbX36+JkWMXpeXPipwTJ3peyrnfJgo5Jgt+w33XhNL8c1MbVL2uaBbKNc4
/DILZMtDzC/RguQn73dcDyNFpGoOe8IpZXwiEpZrvK2Y6KzPTnYmTPpryhkusYTnjy/vjjcnQKVt
OWknP1D1rlaqBEtUkTkFMXbWaeZkS14cXFPEGz/4s74XWpVyt/slzMjho1tNRReL9aKWtlpl+vog
hgefvJeNFJp4xcx18plHq1ey7J7gjvbZuJDs9bMaQGGYAJHc0K79Gpq45Nv9+psxLec1FYKt4FZc
upumr3vsDHd3nqPGeMteRYMYmqoPTxWT/kSr2Pblkmngp4EZcwZsWXCjzNtIOE+9yglW1L0Q9SqY
SjLAKWLTIW8S/qRpPPLXTVDXmv+LTwWQCB/LnOT8qze7xO1a45P51UHqzD4i0h2Z3Hl2VJF8aXFa
xPLSITYfrOgLGjdlLxq+K5UeLsncSDBkS3qkjTy7GQRnMaYmOBZGQSa6MxJfo/mmyz9uASw61060
DrjMaErTSGDK+T/M4EjtL21pTxFUjlSAoukcmtq2tJrCtX6JgMzXgBq7qZX+RIJJLJivb0omdT3B
HNTp9owS4uyzDgWr34sdqCqgsuUzyQZpkbCQ9PXgp0SYrmuXvbHPQWpwYK50emLP8LJaXBrZ6i0t
7UvqKVbVlFawG0j1fariO4cPj8xWUUWm6UYS9FNNZSrprD3nwgno/R6XhTynk5pH+ebydXJNKPHx
pv3LS9h0oRaHeYMiCS39qpOfXfI8yCsA5CUf5GansXLflDaaIdMgiXLx8+dHIsRz4MygPDIqExQT
z/rzf7psn3QTX2WOL7rL7E4eJx0l9r97NBhCVUlVZAric538b4YWwwd8pstEB8IwAVGrE75FBOZ6
VOl6WcqkcL1CC3ok7hVxCD55tWYpudgEoSTVhkR01WeliTllsx7ORn+4l+TzhuVQ3w+lifS362Y/
WHwDRyGlTMftnGVXuJrJLIQpP+dY5k5rs/l47bhEWU7UVIfiPZ5Ohxpg2cOPOXKI/CSipDiL6BMj
6WvJv7ngMXOnBQYYYxWx0sroT0IHl9ZwJcsmhxTWOOy+pKdm8LQU6I/BvPKIUIQcuKGcDao80SQe
4Z/sdIeFbQ+H+F+3dOqUwIh4jjMEfgGpU8cf0T1MCZ3T2bp3pzzpEMZJElFkB/nDfz1jqi4idvda
GtCjkwr9hI9dIAyAshkF/z446NjHn4Nl73QmyqRmdJY/+7CB2G0NmonZ2BQbgP1eQ/GAxfRwO2M/
h4a32jqLZ7wYvKtwyb0/POGd6hnDEnhQqacSg5ZWbcjnxVbQ4gKNceLp+WF6Pspixh3x26bqjN37
qywVqKu5SXNQGycuMM3vHFilZdhhz21+uXRi5ujkPMsBeL/X1VKlbudUcTaZfB2OjF5l/EKmhnkz
JNBMKixr7UVjeSoxCvu+Ji6rUEmy+XgfyR9dIWBjFVH5kUgxVS0tSbzjYI738HUTWi+SeHiMx3u8
izkrrR7xBJAkJtWvfWWyN/ytBt4wwWcqURgQxU7ms8CGEvcz0NZOZu4PrTRwk47QSTwfiGUBuiv1
SJHrtKN18pctg64Jme6xCA0nhQYzgeMXnjXieUcH3neINAnNZ8epEBC37jqI3HlIZnJ1Eo3TgfFq
0gng2r3xILkJpDRJFpmhzJTc00SvROS/UdekEePEv5oNxHHlgiJEXINgBytVw1KpYUaiMBzlRSQ+
U36Ksg6QLkiHPsXXsNYUJLMdrS2rrw/H9UNTj4eIHw8Q8asyzWRS6bvNOHPm07ihyGwmtRcGEh6M
8FHKs0bK83PkZ2IMYlWg0OxImh6ht1Td3kV2HPLkWxicu87JRKKQxtj5tDqXHG4ZoJf2uNu/2wrV
4L0kzBBWaIB2xfShdkt7toXMuoc4khIPbPUq0RRMMKv+TANMINSLhJzSpdg8zt6OpbYoJXbVSQ6s
5rzDGV5Xq4yrG/kwc8SmoCZy+Mfc/nnBx0flU064zNWNYNg0U/qG6EVoz6uElGFSsdEwyjNmsv48
NGAR4MoDbQ17NRVt5fQw+iglWF81Q8DfRdYQKXqgYZ804Vq72zjqBoenS1phNKeslneUZy5iu4eA
uZPpj3sTaG9KGZR0Q0EIIIYnevfAoejuLCMIurptASk9cIbxZ45Lxdc7/rdBRgMZk/iQ13Y2qKWq
gj7WqE5HZvc4/e07vvXGWjf8daCS94LkFUpda9FvBP3w4A9VTaglLspYVrvz75A7hVOz76t8HJT4
r9RtFrSoUIRFruPvw/g8oNuLrDIHtxv/UeNinj9hxexwpH/4HzUFhzCAKq6CJxk9mvSRQ8v54F3f
AubemSWSJDtxbmexKhMzLi4+gMsdGGTGx4R+ijwwKba/LfMy+XbEjUSuesfJ7Ijblw/3h5rxhJGW
FOMTRFa19qvFnaDOoesNdV5qOEF83hAhW9Bs5poYD8RbIvd6sTq+LDjxuY8K7KfOccTxjZuq37aj
3+S+XYvrYXje5pbiGbbfkWZCG3jJNNcMig3BPHCDvvQXoy+9gU4oGn4I2CARz1aSLdymdH649cid
RxIEbmFJKPX1CjLjmXrD3OcjrmezjBSmQSll/7k69wZuUfC+JJ5RGW8fhGfSHiZCeYXVT2wS49Cy
S/S/1wDdAQhmrcefUQKI5rdaO7miiXpuT3ieJg1g+gt0s+GebDJ+XTjMcQirkOca/SWt4wz9vR0Z
9d1SEyhiWoi7Jwgp3baXYUJYVp0Prhcaw+audYlBqRDaaWXZKCC3c3DGlvMUkVXrilFNJv+u9ZYh
9sfJ4ZqyOMAp1EL5CgDi2+vMTJBKlZLiB1TNinIvrfvVn6SZTdfLxOz6IAC2w80n6Im4ESkmmV04
GIY0rLoErfdWYHtp5P15YltS8r4YV8V0A69wioAFr2UZDZneKw9TWKMgqMjYE210f30pgv5vcEGs
CxmwZxRyBCZJDM254aXmCHyQTLvE2jgMuDBbnS9MzXEOO5WyEppn0/3rlt+Sm+qGIt9sgDpQYG3h
lueH1F1ehVL/ZOt5oHMiJbaOczCI6zbqL8MxMe2NPAA/cyuB/yWmcQwteIgyEp/2gRuWAQZ/z90Y
lsrTOF4c5c0Jot56RyOeuJU5RH8QldZAXcZfqQ8iwTVe82TkH0CQeUsEzi+PKMQRJxfzhOUCliDU
5App4EzhMwKdQt2sHZiT5rirmuyM+ov/rQ86tPKNxVcEAsodzJdnHch0ZeWrmGBbL5/fLDxVlLmx
mYPuKuEEW42Di5P3EgL9RVrUfH2E2WPXzMNDMWmCqq0Ju2HAIxEpICDupt/u5yWJvAaj8wd5f8rV
rcqxA9p88OWAidSHbfAwP8ELv2hsVN33otcHdjkR/LzhWcCrxfFBmv0csvVEIsFzF2kX/sT6XO1R
MbPSbvwKJSUi8hwKklS+UE/xCzoj0tGFUSIwy1PLjYUnfVfLb/Xt6mQ2BhsOdjRtnA2qJMu/hinZ
4MajohlmERJyq2K/sCLq/VNrsZTgbmpZBa767xB5DWXQOhiDFea0WU1C4CkaARW7qAL98TWEhstf
El3siw1BH4tlghjdRoeC7s2PTyaMddSNPHnID+jWX0NdfrD8PuB9h5B5NIhk3dRaqeEVOML/ulih
TZVr0ckZz/FC3UIy+ClZvSviNtKLKW+Yy7o7bvAyrtRrLWEkViiO/Mw5cVtw3xJNVDYyGyheqDTk
e4qY7HLFNbMVys8bxOOTgeTPNu+Y2FtN5iiQ9du2cHke+Dvq0BIbyorqbp4RHyuDQeK7hNO/Lj6K
62HIExZ7rEym1ctIds+pt7c3k1d5nLC8r63ELIs3xAqZpA9QGZSu0MZHnRnxGz1tGRWo5y1J37AD
+eAkC19mhZvF0JKGGnKASpVx1/Os0W3HYRfiIfV1ZDj7+Oli9vA1BneQRPLQjh/qtmVUvqj9n36f
KMUYUy+JNuupeXjMmCNZ5f+KD9W7DuAmX60j/0HW5KCBnRw6OsEIUKrvlVvbJjH+tgJJ+kx0UtJZ
kb4H5agrM3aTiF7+88+x0UOL1p7bt8kipL7rVO8dBWYYSgiX/TaOa5i8sYQqu24H4Dtn+YBoqA4V
GaROrld/fQsMO+3bjd0j89o1Q+reIRNByksdUo0uZsdlMlrh/rTHnyVdzewPwgmO+4jP4F8yuubx
yD20cGNYV4mW0AkYFLiVU1Ew4N0DQFh8X7SYMNr5RGUBPgFIBWD79dcxhZvRLFR86Ihc3tT2ykTy
KQ664DPX7q9sonOgkpuJokA8X9P5//5L5TRmtsVPCXIZgKJYxa2214TtCZHMWHCNQKNEdcT/zE+v
KHdtzePcF2xQSl5PkzRdSbeSQdoVNXODNMDPAWxatqOsqGp2iowiYHls39wGnNmswwWW/sOMWecW
wABtp/TlBCSow6RK8xCKdCa8vmpKtl2WVuHXHH9zU5R6HDpfme4/c3taEWoGrgSKX5KGIRN3reLN
ND0YJqPz92gVrfGPryP2R90zp7UbW57KwTGwyOoNS/2tWqJITH+Mp2RoZh0g4IwyO0zjpw4bvUVN
ceDrDKxFBmNKevn+5N4uvQuAQvoGuntzs/UrAgEsCXTXUYHPrszYWFiATd8XCxFPJmBkpFEiRpHc
yCGBx1wib/Rlsl/o1yUKEF9Ibi6Qkme80FLBC0j1N1cSCVNjXFURgbk97aNe6KuaPvWvE+KPU2sy
vKVXpP7Lh6UIGMyQNp6md4pEwUv0on7qj4wSTRJF2z+79QCu0heduMq4vO5Z4qvutZCDRPDQsgsw
2LN05+3O8UQMww971z6O6d7bt+d35Y/CtkfekgMiv5dDjQr1PwFxjOzgfd6jG5j7PDce21P+xDZ3
JcTGtM5Ln1rnKn2CEVPTm3AxWG0jnj1csW5EaoH/YyYF2o/INcdngDd9iCZ1JgslJ6nuSMNdiz/a
Vyb/R8VC+Hn8jZMiqGJiW2QxZrdnUrLNukAKzfJtcc4AneabEQOWyCvbnDmhyQBgzKjNP7F1lT6I
GO0q27xvcNtg8ArCv06ztGZPJ3Tl3Kims2gRlmY2fup9lEqMD3pAt1JZCQYE/Zi5ASSmvDmwY1Cm
oIjVeDiBtWiFIO6Fo9HCUhBUhkYjXW31g9wq9hy6SSwmEz2tqnnXeJXBEh628w35X9R8NHW9kbE2
DvH29701yAg0Sk7cO/hCc2cYkvYujN5WQmJCSrCgqkp+mPWYg1L9q1L+yMk2dfi1k4YWyOxIoVmV
MrCRz7bQz0+FjbYlOefUu6Nf0ZVmwm8iRLxptaOp5838csWLjuohxCRTxVq1eDUrzppBLDlcT7UM
cX1C7W2Fae4HyPFT3pniew3Fq8DX+67RwH4zacsBY/hVMXaytS58QJYi4dBimi4OIWJ+yFYRdQ9w
8XBD64eev8L26Bn5zIb24EAt9YCALHUdPIYVLpECp5jx5ZFRPBQmRL2Yd8R0Me+gUpKbwsBb93Vw
t5DqTrSS+h8e63d+roaPoLdHGLKrzRNCaXZ/jBv9LfHt9/hBOWB7s62Ma/YG+ISKa15Y2LQsZOLO
2TTjGADlW6AOoK7Fi2ZGP+h2ARI+0bzRy8IepvnH4ZIgKIqLDc/m2Bphyve++hSBBmdL4qo8Ccul
QatKueF1IbtyqZ8NldgM4/R+HAgQEjOuD1wtgWNhSVIH1a/1cJCx2x+7TriPJkAQNJx/62xpb4m4
cnTTt+npBNS+nONiciGryjVIPx5MM0SLtyHmh3873Jw/QxOknaqmX6o+4bpINt+eiMOAu372Clp5
1ezr+gP9foq4dJgFRxMah8ZxaxRnsfsD9ZKyCeQtfhEAHVFNdi+zWwMKYIclVI4GmakEsPm2Kc5k
LCkmfd3SdGmxkGTHsGiktpj/gbIC2WV2S7D17pGPIw4yOgXS4RlUKUedbPo2CgvOm2D+nbzfZWUZ
k6dmIpJr1XOMogCqz51mi8WlZE9tavuJ2t612x7R/uWc6vZ8EzJjWH8Inb3ONeZRxoh034a3LVFC
50un3nYCeK7ZWnCkUiwx+/V74DOWy584DmebNL1SEvFVi3MKMM3+UBz39kbEfKxyv7VZqFfjcgPe
oO7RtdYhMMpPZVnhaKqaG0JdQAJRx9H9/BsOk1tEO+NMDYl7CAK5guU0KEmE8FcgpTfs2r13NJNY
YinPClefzDeGyz2uFSjKaGDkLgXiYkmXOX+7gOMZUUh7BTwzxrj7iaJgSc5Vr2l6k8i6+h4+6FoA
hCg5PWYx0pI52KG28MQALUBPtqY6QFeNjTwzl8efyNG2CvvEHKvHGpuCYtMzeuUiBdZzbioH5Xth
Y767/Y82MtPlMyxQjcZF1+ojArWFpCzgL1/T4BedF7mzmcYyh8z5rUECCI76SA3snBJJUGEu3dOR
5PwFuL4xtycGxR4eRLc/18ztnrAoEvW6sF3WTcMfHGOMeS0g7JOPoPehs3ZNvTaFaKeXT+EvjNx6
aY2Z1lEd+i61Q2R7nrTbLVjxUslO4JeBFq3qNn4m2F4BwVq7fxze9Fnx8vGF0yZlSye4ngNcBPhm
o6ahXTSwn4bOW73nVQu2TYFN+FfGy7RSSpQ/bzzp7gVSQ7pm4K60qcgDaEuWIRMZBN9D4Fj5gf0+
MKhMaCrB/049CvZ/2gvrdmCxRInSnA5YfK4HdGriZleSY1nw51AV5l714CfIBxemIM6K7cTdpa70
BZ4i5763brjTPADVY9W5tyb0NeTxBX8k9VWYKvLTDOPlscq9jNXSPoKJkxGBk/zx36b+hZU9tHKE
Xf+VxG1/5cu561AKXOlF5jB+yNosVlZt//yPsGhE73FGS8CxjYmT7Asa5g/XhRpCn+ETIdABKRib
+bd2HdTWMTG9D9s1FR/w6ePYeVSUy0Ey2LGbF/2dEm43uUb1WsWKyx1DGKhMsNDgTs8SkMTfaKPq
wjXb0eaGqRvQyMBilV+cNwMd8pG5JYutHkdl7nvoGGOeEg2cHl5kJ7vJTaoCCsGCaaLosCwN6PUp
uuwWQ//W1E7pK+s1SHO7hRwvMg3l55kgXHIXGkyxfD4iLY2JKFzXpmO7uKX2wRhMbMoFxgkGtu3D
BCZaNSRrxw/VNecOIi600uAsZ8iQUk2xXao1t46WGyFrkGG+ivQw6+jPn+NpIPXHxIfWoCA6Q+4x
Gz+O+NYXkFnchgQgRFV8ESWk2TlsQsOhY/HNpaV8GdR9fs0eCPJD9iyaVwHWFBGaff4pjFA5MTAw
Cf6yeoqOtyAQa0ZqHTx74RPz0MYAw1AuyoPLiNwze69V/3soopUeFe3rEHLBqETf78U+04IxTcVN
ERoASRb0V2Rhb9KWMgIWSsmXDU0Vaey9idH5CLgUgTW2cqw04PDKqhg0dGK0QW3a5sujKhiNNJZp
R4oicDYUhowdFSxYPyT7qX/QpFTQaL9wU5wH0UvThrFmUXX7vyuwxcbqp5+dILNV+cm+n7BS74ii
kJahbU/CnxhXcRBXMkN7qBtgJeb2+AEqYHMPx0BGAC3SRMSfCYUiAAQ48UlgwybEAfBRGd6hf1gi
T/WudJXGlUc0Py0Hh7cKxHYE8TeilNhHZOCUmdyxpYoWf8KxmUT6XieL0/K6RgWjB6eNZDiCN5Ee
c16SP4dIe4DIRpk9lcYG8JEXEF64hjoqpjdYDnQDAK9v/MDA0uhBr72YMckzjekC6GM0bHmve5cr
KHVVxrwknhVGn6irY/TdFrVpWuOwb1oOKwXGU9Rqf2vYKk6cGiZ2hpDPENTTbWXSRVFUfrSnqAI/
tnO29oFef9j9OErWvmLeoI8KgM6RIu+lo1hE5Dqrl+dEU3+GUs4irPuT77oU/JNEG/feUK4Ohmdf
+db5+2s1sIkndEzStZRJQSb40TMNfRHmhIYJVcXN2aHM844LMn+hMLqARgwVen8ghZYS+ymccXt1
Ow4DOyzTraNKXvSC0KyOPAXVOnMvOUPNpK5tmcgjHFXh9tPvUk9rQkWGXXyMyXS+QDbUQbSIMwbp
siKHPL0CIE3sYMqWwUwrw9kD3u3MjNJes1gOKbA8npi3JbpqCYSG9dKnYskAXDQ9R0ddyAcZ+VC0
CrP4P7I3Y+1bEkNkkEQiVmj4btAne2DbJafaiHtOvwqHruXwCrryaNmuOq/3X014d5v+VJbWnXba
q8S6etziJ24c6vZTJr7+9Mma8zOgwwlNTYOGQtntWlGBtGsCx0ZVDHg5zDdv5fTUYxqwTmNbY/hV
iHydLAVrG/Gq1OS5PHX5Gjpd48R/Ykr0rllmh2aFnoQ0vivsZxip2nMU6f9Nsg09xPzXqaZXXOKS
LbVHGHH7kRE5W0ZMI375Wm3TZG+Di05wEP4JPnWcEV46bjs5OCJNEYxkH1PiKZgau/khUpmw0NK2
2OWdnMVumdxWZ0VGLOYXX9tsb1MPI2mmFrDEJHmqOSKGyXTvjo1OaRMqEAykxhrmY2ECjH9Nhky2
uJx+FwpFGZ33FtwBeNc4UJDl6oUk3h7m2s0tjkvMQgOptPhPaAu4lmQvtVskwYPfbKwQ7jNZqUfg
pJ0ItBDeAoOIcFCXhbrN4t9FujzhkvjqdBdP7hbAT+vvIkejS1uDotpezk0dBP9ZOfushrTZxWuS
vcW1q7sjwu4arhb8qQYpwAZhagbMjM9Cdsq2C6kYcISPyCTQbn8SQ4T6fgqN1RuhCotG1nVe2GYZ
3SZGKnwmhOKcndRfU9Zq4JyYneN1Bm4IANf6VPWplxLeh8wyspk9M9TL/an86rgTYnRa456UmRPR
PZBZ6f1EUk/ao/6WwwBpnlxOWgzKVW3hEhnlI12OneBiELPtMhsLeD55x5WkCtv/y2zGOCAQlFUv
ZkCLVkicqTGVrx4ddd26dRftUpm/BU2xYTlURmIl4S8wuNtxiEsiNZXd8PLC/O/fDlui5Tgfzy9Q
3UmA8uyjTqA+wiJFyXQGLo33uMFGtl7eCK9BYqfGcaWwY6dV0TR5kk7Htqmao1j2JHBGHbnuhbj9
fgdZN8CFn6aAUC1ip8tmku0YMitCCM1wZ5Y/COdMn68rDkjGwVZNpNj2NTO+zHJzaWG3AXyundBt
T5DEWLtaGHGMHsBtwJr/OjHcGPR24SMNxv1ezEgVuvFBQJae43MxMkSIIJkzGIoBKJyvD/VZAXdI
pnMGchMz9871olmB04izdOOJUSXSHnzgOgi6nZ/ie0VZ+p4zXDtXua0dRQtdM4bMnxqdsDeEUuB/
MqPYjikuTtdBpp70JTrkd0eU0Gic9TaiRfQtfCGKG0zVI1sau4QFl9czXURfMbGEnTMHNiWZOlmB
Ju7/rE6XRRTYhIWs/c5LLrfp8XhW4RXWL2Y/u1k0b6xEK+4Jh6v9Fvsa+7KqE9afnjM8k0y/6YwI
dMiW/7mRIkHz9mjGl/HQw3SpIici9FYC19J+QIujZzGCZ4A1d5O2Uz79HlqlmNM20nBl3Rb2tLQf
jck9SGYIYgtIrt51wPVTj3LUQewqWLhAyy3jjJjFWDts/SlDkXocJpXX/Cto3t+Mc8jXM4HkuHn/
ML46PDe2wu9qY6uRf4pFPwNVTenAmY0b2022CJNVGo64wcmbMZEtAYlNdzm02+SBvurZ+ithWaGC
S10jloVZSH3RLMDkU+8PUDwAiXx1twIr4M5Y+wcyTyjLC35G91HdnMa3Fbf1rCeoZOmSHWXFfDov
RTYixlrqBPM4g8TeyNOgNy12y2MxHHBtrXJVzutyoSHjFMSSEvm+TTwRLXy7QoGy8+4O9fA3Aqc0
MCuf8ST+ca0iN9tnCmcHqcRtKmLcUqCFWRWHqvu1tQiqf/KuVTczE0RPzyzbxIpoZDpGxqhUyS0J
gZ4GqWxyc5SuBPFbKC7e/0NqgVgQH4iS601gVEmkuoPOo0ztD1UYMJvuTmQefpb2QY0YNXkZqySF
9hxGzIiD+ClyOQ+I2s5KDzFwj8IN1b9kA4tj+rfBoqijTMCJzCgenCYeHRA+erLLtY3NgqCX5Mtg
+GkNqQ5gOXrsVNpdQnp10U4xbnxAwOD/o9VSkchZie3WSHJEo/LLI4KVJ+5nl9PvJljgKSJibqC+
NNXk8zu4M0lc7RRnyQ+R4qVk7auFL5jyR0h1183kjqsfMT9cp0mIC8pIx3YitFjfSgralSUgekmP
Far2gGndYQtJwA0nJH3vC1MfBzfJyCITRkdg2S1fAQUQdKIaqv8zzEP+qi7aBwtren1AyoTO7HG4
YTye4jX86wlUblSc+bUTqanO/zJoCiHq/37OpwgbUYYmdedJ56pPVGDy5+K54gZK6j9j34Gmysht
NNp/iIt3NFbFMqik+IefLaWwpgRGy7DtHEAW7tY9URIh8uw/k/bTnwbOtMiPtB2Pbklg9rTrdGx5
93fwtgjRNUyIfgixUSH7YLdt8B6HHpIqze80l2c0BJV8bDfGn9WqyGlYdFa5JBZdk11UX7W8DeUl
N6b2UZlMxY/0pOjaWG36uW10E8GIHFVkyLz8vjCyaOVC2FzE1tbpKapCm3YfCup8VfkZa+aw13Oo
wQyFnotpIOVtGfJv2C+xjH1Pc+ksm67VhI+RZr7RCZVkTuKDfDXzGyPjH8JO+rejRJy42tk4yl4B
pW3Ut8kqol+7zHVtwv5U3GakPLfVOVdh2zb8S3GlXcYaqocOeEqIILFp+/kHKIpmN7I4gnW47+qA
sEMcRNC5//8CbRKisK3Sms6zsumERnoIhVIOvZBg+qgaG//tsOy267iJCI0vTGsD78sqGDHBt18W
hiOyKvFDgvJYejJYkGTANjHxU+0NtDPpKUdc7yS7GY0XhVtW61baOrAHSLF8WnpKAM38SLeUAfda
8EcTZzHXdzssw0AGSyE7ObWrGMZ4qp37PTfDDb/ml0SeStwc2RQd32xKjkBr1OBB53nNMpNNKKje
tGZNFOgxVlLDRvSmFRs6WQ71rKbLanRYUGy2ZyRs1HVAxdYPRaup//c+bLEoTSwEiGfugVdEx7jx
ZV1HaUbFJDgsUAja3LeP33ZfF100g7gdznIad9tfstjFFzdB8Z3QMRMhL1PkLa42mK5b3Te107lQ
W0GxeirLxQ4SG2QpFfcTBpM1aRCWjLWxO58018kl6G0iCv98o5pOzR2LEtK6/kEyN7fZaNoq9Bm9
4adJmKf29Vsjag0csDHvxixae7ExaUOBXbvWQeRk3wuQ7GsMdGXiD+Py2zzwu8n86wdE+e2OJT5/
2+YPCU/Tq6Rzq2cFojmx837sm0VW5BKFGlyIAGjBWKwO9ZfP7F+qBrZI2XDa9PO6y42V+cUmMe5Y
qghZjlC9BIhkD4nGWf2dTm+8GUMVDDxVmsch9NSzcqCJCwMDRUVCYFMyuJn/Kky4N0Ag94gl8Wa2
Esf85OrwHNsfX2bIOtgpFxtiw7TzRfijIdX5jGIgvBu/Z1hIDW2uPAkcqhmS2+8eJ8Va3XuPtJeH
O+WydVtZQ+s1mYv84fRx2uJGUMH1CndilPim/L+90taqXUK+6ETb4lCyA8+9WMIlsCphgegT6R6l
QX6jckLz5aQV/6gORoxCrlUrMU3bY76SnWwbUKL9v1Oy9ou/GplERy6W0+TSZyDefdye360lRUuS
fIaLBRNFT9H8wDvs/14iXlBbOSoODNcoKF13GHmbjWOQ+Jb2vgRdxOBl+EL42a0rpid2laAs/CBt
Xi+t6F3SV2/71oBjILwgFbkDa5OFlfHB/+/X09kAgs9+B8Z4xGd6ZRUVoK7U22q/+8DQ/br9t8GU
uCQ7jWlxC9uywekOL8F6Mu5nov3i4e9RYauYc7T1DgiFC10UU+lDbVdV/aC0Tl+YlT6szsAAS+8B
B9mwzLLnNIeS9y78/mY3R53IyDpiPQz5MEiOIgz1PHfSS4ns5JlS8IifWsAACEGpO5E4lFrmc09a
Rg48PDrZVmnJ11JdK3tdk5wvnI28Y23gFunDSKkloK/9lqwIy+4GhjOVpwbf3LUfy7oAXUXP0yf/
Y/ben0204AwMZlYiIAVCfXZydHIo8bJTcqnoQgOYCq5NTYEiyHbkIw5T0q0Xag9QDtUEPGzy+g+7
4SCmiCQZvcS/zDjr2olhwcQF0HrZ0yq4W0bdAs2hoiM3UEu4kQqVRJ7/ltXKk+DsjJq5yC/F67HF
SbQkWslpbIAiQkNLYUNUAlRJXAgojz4ZGuXblqX3oTLG3qpKj3AnjxV/4DDK48Bq+Ih+ZLcryzxH
JHkALtHi5Y/NjrqXJtoVueD+QA1U0NbylvqdlnLp29WWBcaFPrMCX7ITCeuY86lNRuQUCk+r+PQw
lyAH31UYfUiIAXKaSRISmBP6Ucls8MRBYMDSPR/Lck7PSXWWsjtoSFfLvkxC1xjn/i8KZXomqi5X
E4FtKTsQzX/iCyVTuDQFDnIyZtjQAfYWNJC8mG0h86VMafZSg0r9sLNc0IIL7dJbAu6Z/1/s4ZKS
0pmPuhppuBGJJXE/O3vV0eueUxNYb0Y8dfBmgWAXDMXcmRJzCrNF5ZqxVzu87DepYISiLEnMpiWu
3WsbE7W4GJPdP1vNMwJYIA7GnIzTb8KEjyn/lQ38fPJs3wPBOzHOzu50TCPrthvgan4CWN+X8hTN
HZvz9PcQ4LuWNnSyuXpr4L1ZOpXCslydwoj3FITVTgX23l1I7qj6sGQOKzpGaJkFPlpt3PId6Z2g
wc+HL+8lFKHwBb8LtDZc+SOpAFnc6JiqN1xy8NglKBMynNGoyDmOoz3LRM/HkWGiy/7ufQD+9f8z
3fw0aTbITBQmzWONVgypIQcw6BzIZ/JJJH7juLa2EsqOpw8MaJVEndAh61q2PbO7T7hovbNgJuSJ
iVRtbxgKdq3rLalSiaYzkJaRpQ0bJbbtFO2PT7VJwpWLgSsWcArN3Bmdm6g+6wqmkTFi5dd+vGSV
CBnk8Q54oYyZHko4lAWlIvgaMrhssDs4zyalZeqph/aRiQuCOLgsCKJx/g1JQvEKMEIHPHQaiJcl
+N8eJNIFE6W+6yNL7lybyj18fDeZK+iAdojpVCbMEslnCJWAIFRe9L2YrezB/8BDMPbqwyzrSUk1
zOc/9QznjLUvONSixelU/y+W2B36XZqa1baINoi1ejea0BzANjLyYfwPjWyTHxU+o3CeRhQXwIFC
5g47Q5m/gxht1q2Tn9CjtSO0qL5HgTYmSBZBRrpo5oMF1imfJHguTRL26jrvtt+eWIGB+90Opso9
8ggP7T6xCyXpUhwd9/ef/PcQeNWyzV1gLP2JlyqPGNycsS4pihJuOV0H5ps3VZPQkD7q7/oeUSqK
kLJs8QIBI3A7dFY8cEaTClEN0Zad4pAs4jK5X1cr7zna12rfb+hw49LOtDvljM5VXLeGfj2y8ay4
4a3FAEqUmVP41L7XGh5Xm5fC8G2hHoMbCTnabYBjCnCC8KfU4/LDls6U/RZNifMYOFZOjCX5o2jM
pwk8PiIYpZINqYP9LvrU59lqPs8Rip7NeK1wcDaDuqAkBME/m+XYrk3+h2vrr6ZWRI3pu17iJKfq
74zjT5KADSvHFGvuTYI8t5jD9M+sXYoyCaJswjRHKbvfTXyL9Afdx3PjrNhJ1gBqLHg7pTD9rYCD
BmPSn2gbMZUVbm7i3cGxR+MsjsxvF5wA7gGryyDdmvLLXmrfbOkuF9VAnfFwL4PkYCXQnIEtZd0F
LvOAhXHrACC2OvonYnLGjGJH7gaJN9bKdotPJq9kPs0wvfbYlkzszMP8+aTwlv0smpP3jSTqkWFJ
PnopMczOGONHgZ2PQQUg9UtUTyDJnOdjejKAEWVZqi5z6sb8rR8yX2JkhSu5oNKAwyh1VvSTaE5p
TD4bhCk2fZGZz8LFZbAPjY62F7gvbeOSRaLRFctJVcAXUqNhet1P6YNOOJxNof36PIh/rKd0+yyB
6UGFgzyvRj9YfezL3zPnFqdZLQQ+LhTNTzHsGmL7dsoOhCswjrfEgODC/EWn+DKRL3KetwdWxSO6
6nsVD6hYeqjnMUryjB8vAQWIMNrOJrC+PCvvcKGJukA7ZJVmtlp6UArfo8EpvC0X5G+6DHT+2JFO
KZqSiZepvucf0Qy8yBybTUIWT51xSpgTOH3AasURsEc6Un2sP9+qAVvHOsBlnD3N8r0yo9//Jv0Q
5hkSj6QsNM0cY2r9bPojUh3NNrbA3HPPNmgYBO8yOqjG82CClVFDXeqzEkDIvkFQUaECe72GERGC
4n7KcumnJHdW7NT2RcvbAn46bAkbJ3iGOi+9IRT55m1ZnHKjG4d1lKqFU2wJ3kjZRo0+yBrFcEiz
wXGqoPHRj/p+vUFzBPA5g+SE8R1Gx8+IMJMmJnxlFQU2usmnKFgtHBSykTs0OnqI2UqG/k2A9bNz
fcdQxw/HIbpdY5FqwqqQvM9qiZwvF1Ey3ZqYXHiJj1nw9mG4kBztWsDjsOgzYSLPatZ9sqYKxYZx
qX4s+XD007z0tI+CjOkxOVqfDMRefj+CeYxX4JMvu7hrZtI1lf/UP6WwEKnjFUDKdYw/DezpiwZL
mN5bfjars72I6aJ37V/tDJIeZDkxogZ4f2oPvAo4QDuqIc2+wrZ8Zy2NwqDqQ2TbJsaUTg5SrE+W
/yU2ITNft5QhTEKl2SULUUj2tgnc1eTl0XDGPTtPfybygE1sw8kucMMQVoWDlym3J7Cb0YJnP1ZB
cCwP1RXKg9JB/NIZFMHMc+pHPSzG8hVb5ftAN08Nu1DWB2gCTHALSzka02/5HfeUPq/V5dBA7w61
QC0oI6OiU4J9hB8FLmTZEdwrP/sHeThygCeSMcPGxoriRbsoAsavzMQhbJqbK/MYW6EqOQUtYHAx
fV6KcVe/rKI4CweRbgJSXQm8qXhAyZp2A1hIs7wF1pHDa/y6h0v8ATWo9TNa133MP2WXvNDQvRTA
c66cJekSqAbBDlgRCIb2ApLVGtPKW3O0PiHzoc+XBigh9HsvXA9BCEHGJWOvB1/rTvaBQ0N+pX2f
6Ul6p5SnFCpP70o6jaZ252o9P/daRpQYyeS31GZBkRufc86hlKe4ZfjuOo4AnVQiV8R8ltavB9Gp
7tXgpaLNkem+RPDmt6Ge1wdFlGiyw4KdBk2Sgy+0MEZhykZpccZsQ5LLT3lF7CG7WA2MbwtlQgNJ
lw2GrQOLp926IOrfC7fqBvJOoFBZsjOMzRnJ/tA0YgodFC1drrXHuqdQ6ncE75oFrI+MyJ1/TFxj
2y0bbMqSu2RBNIO/UautM3YARY2GKC4Vg1f1ODbpJQyJjX2rl4wGIqoRoXIpsUVbrTwbpAcXCJP7
rXQslz3li0Tyd2nAvU0VM/jiOzlABDKIAkpqeFf2/p2CmbVkiA2CdEKjZLZrItV4cNVNkGWCalCU
pyjFzNy6c1v2USVObhIb0bovG6ka8E7Zidm0nsQYWUbp9ssZQsr706GZQ6awDib+N3EBZfCp5B4h
guFCzXhuq1KTuoQ7BjClIGZE1cRQvKvQT2QNJStR8MjASVGmngI3UBChThwfgoUUSfOi2oyTvG/M
WfudIL2skAEsXoCcDvpDRZ5qEFWpOu6YOoA7gIsgTJAubWQ45RDzTrHJsakQj9eB2u3VB+I4WR5a
EnEvZmGaZByvIR945Lgbtq3KDb45Pc9lne0ew7tNmurthpnHeUm4ko6IqEN4uCAkhPCKjnm9m4kO
YoUQ3khxuhLyC3yq/XfrW0ObRjHiMhr47qygISJOsNTN1aXFSPc8EjmbJvAg0wt5KQkxSGtaExAg
eIIAs6XS7eCVZjz9ke0aV4+caZNJSo5BFT5kvXKR13H1uBRMBNPqhP484sMIcvPY46GZOCL92YXv
gl/+09NXbtLMTjJhKujUtjhoTWPL0fe8QJzvsAUvgw/zHM1L1sT1KkpPammQP41ZMvo3KguyOiyK
atehfzQLS+odUwQoNMnr/6MObT+rcziI3a5pdcIGvB3baP13NYGWzu5weMLYAJOWH/H7lMPiupRp
ARgTqiRjy8iiKCsnzunR14xMabgHLEZDqPCCniKXI1C450pMlF5Xpcx1yy7wEuoqb9DKFOhTZDNR
IwMNx0dRtC4gYiFALatg2U+nNMm/fV5Kwiw5xdoQyjb3tZlZzmF99bDsBfCLOjQjEYSkZKvCfcej
widZsClnmMSH8GECOpfKTaNHTWvcHqeHmECBA8CmeyUG+rugt++uZnoVf54p5Z2TTtIi4ssI7lQu
IlMKfBNlTxH7PpkcdMohjkAoA03/mhYWexu2ZCTYt7wak+10pFsP0e47ooRpwYrw49NXasFj0fI6
6NBmCdOXjmoV76siaia/P4D+pjyErNh/q9cEytIcmbkVq2vmMNn+60UE93j5IlMrz2mMRp1zEaOs
+zD51jHF5LIfYILapUw/5x1dd3yKj86e5L7eNGLUZbjKMNO79ZLTISeRvDehma1g6dsrNP+g3nCd
iOvMTYmFOR6kDtvraYkXt7GTaONWX/lxUViTJKYu2aTdkBpslBkgc/u0R5UpLSsJnjwNd9zBAEDs
ptTwvkp253en9moBOnRVRz+uqXtwe2UmENRP8dH0S7Uz6he2CFsIegP65+4dHVg12Zc34zrP784Q
e4d7UicIpOJcKDPiRaAiBHxyPyY9jtt63g2vVbxE9RgpcUNuvEvfpn9XGQSxTJZIOR4yQFbr9Bim
7TKGJ/Rpf2vxBehk3cQT/cCHDTUdrsKEFScGaVV68WuXvuQjqBs/7YyC0V4vPEf9RA6EKEg8Ghru
VITTiX9FsVFzBkQGMlsUO2bo7x3Rci/q+zFJxZwvVlqTCoNNUf9PueyeuOAg3MjZJaAbZi/himv8
RnXAjBraeaMv8OOfTdFv1dw3v8r2EJaq5CxCdqGKJypGRX0WGC0Hl7yhUCr0FOyy9WVDIBAshcIA
L/LAzpYy+RR0LS/INeZ5TvKdwfMDfwepv5+yxilwdHwkr6l7Lfckz0ZtVaQFX1Lh76UTAphPmMWC
8Uj3ynzbGP2S5yzDBsWURywMaBIyEVCxvpTgp+XGDWMKmCTrIm2C9qMsQq0pMLUxS7FYcTrOmzUy
09bKQzrEed6eWwgLMWoqRRhoivhiV8rghXUaCrT0nuePtnsERILyQmeVboG7N5q3zA7jvNIPqAQL
jDC3kwceQd8Xubu1QoVKaAOcQop9pTHTLWNujry4+Km6bAxeOOMXWHQdNGTDtCJ5t6+jFgdwd+vv
c5GQZ26MIBHMslFDNCr8KyguEbXbsLuObhVwAJxUXw9rTthjqDrlp6wQXSULIuQl2U8v7lDtvehe
qgpvB4ipLGt+I8ufuJoF8ILE0LKAXUTXu741fffrKNgHBzEgUOk4lkW8ekUk1bX47IvBen/50Amt
EQG0QyUcH/4PraBizgAJHbuPOcj+YY/t9uK1ptXMaQ+op/5COeTzk5sdVz4O7HMWg8o/7q1rObNC
MAXzdm6Ppjfs3i45zaAdS7vIIyBPVsA3BFOelMh+T63jVXtUWsehLwoXAhKFDP0kcvkA3ptgM7Ag
pO4lW8VFOsLZ0uN80CndqJ4ThlNTQQu0rU/jUQeUe4MoH7noth46cxYj3icc3cpSBlwF3KF2vamx
3UnzpLRdDuHbxkSY9+FOXg6xeZ1i00sGX6obyu8wSbY/OewkJGkZreXxOH7Y1flhfwZCGSF+lnuF
N+/bA1oovg+uMero4b25HXQXpNUgM8G8pAiOyDiHCe0Nlhy0QQjPjU7rmxX7fks579a9iJVdDR5J
ERdyfnVZ0haOYz0iTfCjmhsBGKDooou/2wou4qyoJG5sxUwB/ZHOHZFoY7HIqpEdnA0M7Qy8jXh8
MTxMrcafsNlvB50Ign2g2E7vx0nUAYj6MO5N6MgRMobXKG2WfBZr93RSoCBWY16owElyPBKiA6o+
sD2M/OqynepBwb4X8adhH+E/O/XVgKK7UBib/abqH8TlZY6v1RBl9I2rYQ4lzq9fiRJhRCEK28wA
54bOAF5n740SZVCrcYrvRA385valb3zqihRd24wnMW4z2uCS0zsF7VGz+lwqgv3JapqsaQqrM2GU
slc7U5S3iX262pPFlaAf98bfzMCBjhg7+zHJzNnadBqhc+H/p2/xD5vqzPFpg+9pwCnVBBQyFewR
aK23jcuZjwdPkI/AC3BRSaPxF0mDFtlnG37i+eQafF0sd0udLeA+C/3PzRi5s9oySMSL2qRrkHkb
+SOf9KYLpSGV6lUixu9cC+iwFtFFt7YXewMEvjGl9h2m/MPz+PTueRNE1Cil8ExFFsoafQUhNbXM
k0rnHuwqVFrzAR5JVDJbINGmSOBL6qEa2DOAr+hJcpWihNiYWCG0TUpskj49sBWBmo+6T5n4geUs
cEKFJ5dyqNwH3q7LJtP/fNuzOtgpuO0d3IMaiaOrAleu+lELG+2XQryh08douO8/+qCskekXH5YU
WDTip4cPEU3ZzJ+cIapp39nwO786lZpDA3pXGZqTtlr2p/LezewcxY/u0qmbvl3S6pCMvJQdPI8o
4L0OHolfEURC5+WsdLJ2nVnVZhG9PDIzz2rQSqzaxF0Dt0Nepl4S4/oripxfAEl7xMi6yxZjGfMZ
qzFQwMkAyd/8YKHCGNLaEtQzbbqLetDEj/C/MwFSa3c690+h1W+ogKfY2HVS/5aK69AzemVPbI9j
TGJzs3HWrZY+QmVcbCtq1mkk+JE7hdOfa/0fIjwkcIZdq7QMZpH//xPiADL+zzvHCfmiozOEBQ/G
nYkSk7u4YAPfu+4GvIzZ9MyradLa7dFEUVLAxqVs2zFnO3EID6ZyAYjpxkrzDSZ60jzPEkO+WH0d
TqPBWDBkGas9rMuLfXYIdkZ7BNzn9LPybO6tl0aUYwXy1sjDaTj++zXeQLWo2f3TK9LE3YQEYLAY
wbCeNNbknkBVAqVZfC5RGOL8q87009fCQLMm6GZVmXOL5Y+Ork8SFtGhPfOvCXzS7q+0OmchTr4H
7Yu5YkCKPyHhDkwkEckfqBmayIIvMIVmf6rg6MNpGCiM+2a5McG8UYh5lQftU5LRVtURPoADryDI
xBeiwAYK0W5pWq5yx4dUkmvevnbPKw2aLgzOfvLWlunh8aDOMM1ehSZNGeRUsstwaXUx/iKBOI5h
NNtsUGPH5lJsEt4EJb0ea6yA5FRQy50FB0kFEWnk9PUz6uGBpZ+eQiQwabj6q4PDDUTALcDNDqFX
3SWLilD7+6PXP32JLZJ7O14JrKWVDiVEZjE44YQWnuSjjH4QOCTO1k6QUjzumjlDn3BxddAqpBrj
DLSk59iiznRdZiZnXTOxcl7vhY+YhIGMlortWDChBiS8K/bpwEPJS9ivpXSr7XG4m/1D+PEj1oSE
RNz7abOn2nHbXQuMoeOBzJGTeGEUSRLCjjiGvVCVnY6Razz1w6KvPQ3cm1IhYwod3eBH65bHkGU5
dV7KVjUi44MsSyjUl+frCdS2XCQWiKrF8aIUboYbVcV/RexcnVtXvRd7I6Fe81XPaWXLWYZvMcpe
3hSi9R3efJcf+vS9MWnaCHLHyKS7z/4yqaUOdrgPDnG1YVGapkSbBroG1gLUM/QbOYvRlODJbAFc
ZpqUjU3/UvtxwGTBrZsutrFYqGuy6ifmtHA2D1H7OSnj6U6oSWKB6kHhiNevl+7z6cs1rGsf6u2a
Vd8H5eI3kmC3e44HDHtfJYdBEpI4JnhY7z6sbKYbturl5C0AKg7Q3DWSdnu6fkpgVO/Zp6Xa+zd5
Xkf4Ovjbs6Xr1N4axSjnRZNSzLjFZ0gJSz8cy9aKv//qepafE+FWwh30CoCdoPXvD1/NUj3FwLxy
Wsh23W1tM5HexX7qUPGyJxhecnOUbqvORQuahboktQAkaZriw2Iq5IAcBzrDCwObM6e9USt88+xu
6j0QP6bg4ZtGU8qgMFjbytMgJSA2Kp7Ud9bNBET4mFhntq4pkznjZgScgfm+xGd3YtfNHQuiaXcN
eGM5M1jVwUNq2c8/d+WhkGjWB6DDW6uyi42qQHihrRHV0phmQHTRj7o86UWLluY1yelQfZUYdusS
pLneOmrUK25DO6G4/zfpE1eySh9eX36H8gDgJYgT95KCfsyhH+gu3e5fdc2ZScwgdDNRbd6iSVgT
E8Hrha8t1HKW5UCDKOWf1ptnskZtqAmtwlGdWuyRCcPMt9NxLuPsIIQl99biS0zDPfM/wZ6eBQ08
7YDxmjDejrIhQ3FB+/HJaVmVslHFN5Mg5svwVZPlCtmyAUxp69LaQugDzrRdHsnnSTztHfLOXBlr
P2UbCjjJF5+rWhp7ZaUrLOuZPXp80Jked3OfkOMpOz5VFEY0LNPzQ4YbIfJRiWqGPhuFWbcKdqq5
hg0eT+7ayYSl99i0yYi6az6hyAnknntWxgCAWYvboFL6AnfBx74nVQbJhjpdENvO75hVX3Lb59sN
4M28incoepzKPCyapXvVP4aM//OL6UBOYYOYmvP0u2Ka4HEDPupCbQp8Vv1YOXhRSljIUT0mB3r1
d0jtZC/mD5gX2RUJCMstrmwPuf9RtsPOUF0lkY61R080YR2GGLJvgUJCFv/4oarJ6Zt26E/n87if
IVY/lKKWtHF6Oi4NNffep4pyuOos0RmalV7PF2QmVZ1C09mVe74CrZCM5j0SmVtVCKVd436MUifE
tT7rMrShkju4KC2Y/xTwNyhQrRjF17+qsyxZQAFumL7UDvpJ+dCUpVswwGvejRgD3M8dNH0sEkAG
bOI1RaKYWgyQslUf7Zk/B3DeaAMT1QSRCMjvra6RyVpCBPNcQcXS2mrVZw30pzRKYUyKxrMaJeLY
goVYuZB7YMg1TJVcqFksP2nuaO2NCj/+gtZNhxipN1x6t1sIa+dAyUXVYVZ3Hrk04uGdw+tTximO
vXs7jKs2EEm7w7IJ4Oct/IyQ4EEGrIsDsdqDkYo7xVI7DgHNpm5Knt53vtITLxmcyuAUkPHvUoMV
5rwgf36tmUBqeeZ4wwLLDeoYCJPUY+PRyu7IQ7p1a1VOVFF3ABS6IBXyhflEanZJ28LTSBmt6GxS
Cm83RFoWCFFMI6tzjQ+gx6LGNy2jTV5nr3HnlpiG5LJ/TnCfJvdCBHDddJjEUXvcGF2tNJtDChIx
2kqyni/+pm3TxsxpHwyjEa7pDBPK8ZwCuNX1WkMpSP57536b0Ys4MPNHbpDMn7a+5SpVi4tre7Jh
Bh+iDIr4gs6GbWZCWGX76T8fnDkTxtj5QhWlgoSTfni02Pi0fPW6cw2EHwlB5KRgQ975p9LPnQTR
yv7DAB871HmUVCqI6APpRvi+n0QGJzAK7R5YGpk2WIDEYHwAoa6r51WesoWrlmOcWfGi4UPDf+Rv
tP4cp2L8aWd9hXAGPHJDJHodTCFJQGaNUelxJ5L30zmrC9rUdIAwll295KjElSyEGQbUlEvvPC4w
cdr867/VVT31y3JkT6B3L+T6XLLAWnMFLurdCd+4CO+T5EmDbZcNuGTZY3RBLwiLMDNUiIAwLeTF
z7Ry9HT7awJGc1RHOU5FsMY9SPmcWIzb74kDeuX7i9r+ma4AhuN6YF+gLkNQPX9Mr2M7UjNd8axX
7h/u2jSYGTKW/QWo/6Nx1KUNbBjVOCJpjIT7VGRM89DBXKM+XcdqJWBIt4vQ+mWcIsHkQtd+A2ZE
VgWSj0GZwSEVtGcMwmlupV8ZamQkPBVL7Q2scPBY9la+4lftPziANdHG4vlw4U4zV9h+pREaOKAH
36d8FfsiU7/Blzfhtfteq/B6JihxF59WMmJ50MFHflFX/5IojD7nveWEGDS0rmHRAbGSdvZwT6Zt
DjZ/U0ZSDJ6NJGP1hB6zVdi5y/3cXurM3WfX8PYsxoyVIEcq3AK1jz0R0Z8bqzBeGE07xTiVZEkh
shuAVJAShFVfZTnK5mKE8X5EbHY08CesGi/uCtz5PeXH5VKQdQEVztKknyGrTN2tDR1E8eDm/CIV
bZrY9gTl5Sr6Hh3gQX7qDEFtKzzFpXLxGgWLS/sRHS631nJJX8uVqDvIcBEAyV2Yq9BNeM979HI4
BbLLwk05Bu3b92lxp3jJctFOscG4aqs8QHazqNlrVCiCTENDWqpSeU/eUbIXi0PLgb1uCZAAH+Jh
VzmS/KacTHaZ3jYKYkIFw28pgBbh6234NAR/yOLEn9QS2cXnNdc8WOnx6WsaN7KMh6QfSF33Fwyn
x/TQcSgY3Yo6fyKRZnzRdtD9QBNPYSLKWztqxL5tGLA23QsvGC0XfgpKXqxMxJmdy4bw8TSflhwW
Lxpk9gzsEXLFqc5yLi48YRXBwSi9f6nbeHo97S6ZfEImNwV+UWZ1Beir+XwNMTj3Yv5GT9KrWTJf
H5v6SazT+9EVhO5+FWPV8Bl1C9/cOrzbS+K7LNMzSeAIHgxBK5HvugQ3mzPaLke1GYB0Npk9dU6Y
8u+TDBce5aGJwGnT2QbGX91T7c1aoqO0UjMM2FuHjVH5X65A7m7MxQpFpZltv39S1g29fjt3yho7
gfrwUJ0R/o4GNb4bNPMavUrPX/yWskHgBqGSSPAaQYYXukH1T28zc6vH5T1OAHetlGK1cYLA8Mhh
FgzyXqPt2Jo0vab3FuzzGhgeBy2vShHHuxHFdlEIAxyxe166DI7pYegXYg5ClBg0/GtaPD6oNr36
y0ES4NlWnJOQG8VaZPlByOj4o3h/vEC2HlDBJ3LH7rc5LBVH0AorQ3RVa0Uo17q7rk0+xWB1Q620
n+QxkPgGeSDJG14JsqQZx3sqgL2FKaA8NgTiIVVhHB4dQI810IeLBS0CZVHnypqpAC+xdWSaUMS9
Y++QqEKBpneOFc7SLZfDFvgUKvB0s03JCHOttO+/icUYPfpVGZulm4xT69i7k9/yrH56bc74tp3P
H6WFz4kSq1HFTw+mcBj1mAXr2yOnxkeeMXly0VA5xf8PKDf1pnArDgMzegx9PXDzEYYrPaXBF4B7
PZfR01sd6hpnG6xO8SGS0zM+VFSIGyLX2ZaAxcbivNEMj6PKH2KNvAcHvYOsRVwTpcNjHcCNFq1L
Zllkvl3PLoOddDexiBd+YdVBae7/7Sxu5xDRc5EjfxE765xHK64FTPrrzBbicwlfAdt/62imePCT
HY/X/Z4skN403hxZD6PGqoZKZxtoNyEIyPjHa4z53AJGmZ3JAVhq76K01s1FrUUKe/e2LrY6w3SU
FFenXLIExgI714GbMRmEWq19OKu0nVBrabSvlMOSzO0QBLcH0pNC8uUbBGxfRizAmafwMwyXqSwH
hFs7bDSDPXFx20l1og59T5A6DMn9BZFQ3IPjOtOcAS03V5cPkzLQ0zyxu9C6rIL6xzGkWej9keyy
sI3Y3sSEb2hXhRAdWZz8GASMDsAJtZuU5S2EY8RUwxXoYdt8AjEQ7l2bsgwxbKgOvyTXBzSZMlg6
3jXAlh9/0e2FuonmjDlaMQ85suz9AqyYtsWWNXebogfhINdgU3GtvsuQNxAHewWtyh1Ii8GI9scv
Wq65vijTKRvk4D2df4W8kWEZZta1TvXAGHb4s/9rL3OfcHnCl8+iwDj4dE1jJTOqn9l3SWiy2hC7
ZMvu3bALOQg8+7lXSVZzLq4ZgsXkbuftzAZUgyfFfoCfink0sViYJKJt37GZRa/9m6v/pEy+D1Gb
jYpNY5AAUDAwRawIpHZii9UJPX9Kz7r4IWc2rT8qiX1OkdR0IPChaasksMRGV2C8Wu6DlgB9N1RS
Wx02mRMohQ9PXwwHBUouTq/HhJh2zKBmafhBHD7sWiySTajVSt6wR/AyZjB6eK3xcuMdFOlfOFy5
nShKGITTHm4Q7L2iNpciBP4nL1GsrBxkB3wezc3juWfTDWt/JqRyhITVN0sYT78UKsWZM61HYHAO
HT0A/VOerWEDp0KCbvk2us+AGNc+CGW2JwOaXbiDj8Rt60PrCiA/m9mnv1UBLnhRBAskKiPECYSY
Yg+byiPwNWDWsRKmMFolnPUPlwE6AdqgGb9Ah7/iYntkXBS4pTpc+smk3rzrO2QElvgl+WXMbVxV
7d9z6KYVG5UMzx7+A3Fhs5veNa9tbtBn2Wgqdz3JAqTYce9K01A9uecGBqLUIgEh3BeV5B75HZg2
2ibgCoAccRfnp82dR5ZMtgrIgEpbCU8la+8VDsVlxvSdWJnjtgOJ1igWeYMTTzR6dnqH/bszI3Gz
cqeDUfVqal1rC+Q50Ee6IB2hAJUQNAAtf1JxBJnoRb5YhCiL8rHTVP2p2aRUL3b9lzbOUcRXHPEA
bYk6lySOGmYl5mvsFMiUVL8+6N69kAULkPjGq5E275JM9Rrcf3Tl2e8GwN4uZfHAT3h1BJkzWCN2
KkbToyNbZJRVjLCIi+kq4rnOzrsVVNaTQ1+SDsqPgpiHCCtlnQKebsdyFM5SkGsE5liBjpkcLq0W
nTSlXNPec7G1+G/xMPDxKgakIhD1b5m2asWIM2I55Ss5s36OqD9RWkiT7ojPSf/pmrAf5p8wlhq7
TLcSYiQg+V9m9DJNR3ncNNTGTDfrqvVwqjs0TUNbwELGydvvX8zEfsYz1aVVO8TY9qzbZ0wAhNXd
Q8mas+eyAHWO129vAKSuS7SE14SahJN89C3Sbz9h6OXBkdFbdjydc2QTajAh2G419VBpd2rlGYO6
504nfzwzarw+wdPbQ0dksT21wvgk+2/ChSi1gV1yc1qBYup3daXYuRw/tJocFbhe999ktu6ECKLJ
sITvOiFKfdu6UxSivAdO0pl2QM99BahtasS93VI3ARoLSIlgC0r4i9xgP96tIduRjjw4teH/cI0C
PKo6kr34h5BPfovg9hKV60yOD3OUWmjbyEJ0Y2OJwd7DhY+GspDTwalMmehzZMQLyvDyzPIT2YIC
iLHPS1EElJSEvAg/vinbylFlg2/Y6tZ2DQolxv6NlzEPmAgb8LDawmUeqduCguEVNJnAulkJZWds
9wXeCkUNji3osPKQIb1T9r78hCxz9G4fml+GXvHaqJI+90w3xhwlDL9MeSYNEgrMVgAVatcCq4/N
a7yQR2fwY0zVbqf0onJai4nD6Ovgi5g5uk2TM8uLGX5ULMkPIh+blAmGh4QY1noXtr5Q8ewHbYZF
5hkYAR1YcDBanid5BVdq+49F2agBlnlbRSePJMfRmu6fXU9UYAv4uF1x8ftmwFirWadCluGp/he+
4wJtou0JED6ekuupyxGT5m+G9qU8ZBnM4dWZpaGlf+hzb3CCYzdIj9iJQqMBGRLNuabZjjhBElFk
ktFBPFyRwv2OrJKD5s9iHUdoHXafn0bOAKrtdwwarP0G8mNDeyF9KyTbtF0BoZRYDBzikRjOA8YU
Xw4jgIQJAy5OlzuU37t7LDnZ2zB5AklnKZJtfRuTQEUcr6N8b31yZ+5uLWtksCXdWgKmtPFzHZYS
8sufaJ7ypQKfAZuKF0ouIwh2U/DH5o9daeBCuxWiIgU7KJ1faleaB2JDyMGNMnx9tEUuBu8hQhay
gng7HxyWxO9wHfUdJwO2dyRpaRHFx5KFwe6HyqXLuFriXzrRGs94zjYse3OPiEUcLeIAUQYfmYRk
1TXLMWe2kooE26R/g4b7Vcv5XnM0RjGiJYTK3xZTX+Na2go9/whUZ8zXmGTYM3JcapXgZFcCYjj6
XngYiCf4KUBjKgZK+paL9DCOjy0MnLMgGg81MYzVJolHtLdFwvcCnPldqz8UfssY1A7k8lpKd2/Q
BXZICe73OvZYeZAYgyg7dZKZc+GC1ezzQraKqMg0zJuR6J4gF24RVc+8mnrbYC38NrLt+zkBZvg4
XoZtJytTdpCdr718+yuUP7X3JELr6niy3npuU7IBROyk8fBr4AKw7Q+kxygxOjWqpvJ4t11EcmO4
+ytXJoRsSxtPljtpZsTFAOCpICKX3qp+S/9XdQMJb2tbkkW2Tgit9WSELRZrI4FMG4ZKT7+3OFpM
9tl9HJzTKECAOjCko/RuuQf6cIhLkJLONdmDhfA87dRWhCHI1AB6yWAytSIiRbX2tqBkJ34z3tLS
AeCV45TrtkUhFaMCPnf85rXRkkdHUjErTr+0cQcHbGowuyBXQrg0Ep2L7L5S+Rjl/awdH/NZ1X7m
7aPblLq7IdiKHzhH3CVvT9esgo9CWFBva1LMxcuSdEK2ASdK/B9rv+RzdWpC7E7c+I4AZOWTOXwF
d22B00eghkdSP4JDND+MYy0ZBstMpm1/n6xqyF/1pUAB34R8GrFRwweRqCbeiUVOD+3Yr/8JQUVv
eOk+awPSNxKYqEsp0nyyOVxaVOZbxkijcY/TZeQvUqLomEzbLYjghbbe7taqC4jD68kW76KBt0Zw
gCY7vSmtVkDL2oW6+sWnRC9nMmsYexu45GhcXalVg3vAHBMalFBaWXenzI1xAKdSvtwuOIMvb+Cd
6pyJCDaPla6MZl8o4ctwG464wriUMns9Ab1YTA0PPja0mAcK2C3mzPbwHoVCDuALqAAPBvvc1idg
vQHqkUcPwYN48lkKLkXCiE8qxh/ld8c8EC85SbeY5dsoYWirci9GodrnObyBL1givhgafj4uRFR4
KNR7eR/qEPoB1rKjyPQOD+pZR+FIlUfqIbsS+GUJXThJE4FzKa45O6nDUslx214LXnZ8nUJG1IbM
yuLcRSOxuU18zQEOVxpMEvzMcMUJFnFZx6ojPs9EYBoXFJORK5bDupup8+pGIgKYhdXSqxBjwlwg
6bYmocPwF9UCO8BjSNIA4OIdYfS0tYTQqxO9ImYaQvjoyrbVZcHUqpSz6e1/tl9YukxfX4h2/l/0
KhbC/4xok3XgpU/HNcxB/YGFwaZNbuc4hdw3wtBFDaN+0Dxq4IFBIroGfisYlr4M8gDTlKekCk3J
bnXQy42KjbaxDKd0cP/Yu/IwCmD3KBtEMYR6g8qSS6laWqm//v2DOAgFHrUyq0l9X9IQ3mSzdUIi
aoE6PpQT1pnqcCM160yEsHSOSTUW0VYwG+hUKaw2fHjOTMzsVH94hjW2bE3s9meWguFd/ooFu25k
w8syht5Rss+8Xsqw6dvRoInanUGvVaOfagzCOu7VI8kWLJm/93p65Kh67hhwjRC4/NQH7qAm0v2D
8KUMUpLh/UTg8iOaTBQEdYjb4R7EX1GR4h//XwFlqHmqjGQ4O5vcTIRnhRmVBQTZmYwTsGwmVL7c
kUiH0xabg2aop1GFfkp0HgsDGZ7UGolgHt4eXGpmmDN5Zsc35yqrDdk1OoNFYDIWqZeH4e4mYQGl
MjG8PPEiByaE56VAT1KWLU7kvA/+qN8Bom3MAbEB53Rzt8Sf3NxXdDiRI3s7HXzPOs4og1UO1ICu
QbRAgv+9CUtsCxsRXfneAkD9DtucufKBvGwBEfarM3LZiETBT/ijaTqwCKsP4urzZErYypRwLx2d
I6jVGhS7cQ/gaBiwlbcZXDpFwvKufEhvzXxhc+zNQkT/iaXgHaNnNUTG4nSqyMKxzX8gfPb9euVx
5DYaqul8JejJnWOmoSxVKpjkrfAAhEP+jnSdvW8A2cool395+R9V7QNncudfGeRz36CDAdkrYnvQ
SyCxwbXe7+POnBRJzC5HEvHkX5PVwTwHE2cPGgCwqh2k/LIY1H6sGIobBjCzJ9p6ILIBXIhSeBkT
iQceZ90DmJ5A2pnwIuAi4AhitdfCg0EK87/jeKK2Gkec1wQZpKAoItL3vimLsdTvkzZ9o5LG/JRv
wVK9ue3sjtoIl6QIb4iCv9Z5gVHMHRJCATHjtpZext0sig/+2zYBx/wfgoTs7w5a+mIcP45bBvGn
iknDf6RmwN+d0o2naj9pG4lqv3+XKEJDpY6+iTwknwV5RpZ1JNgz7zemQhZiwuDPHTGRDFXwONYg
EjDHG97jgL7M28lKlJjxTAVh8286m87uVGl3IVjvoVFpGtlUrhzvxYchMqKPeV4d57dhUsVcnM6l
V54v5TiIjHERbUp7BylrkJG2z1AxA6cffllrnlkVYKodtaupDBY6iZwo3BpI2uKeXb4HGhCJiR6v
+gbV6CbDvIXFt2LdHdAW/uO/nhaV43FKAgg98ixQAxw90mOhMZHAo+ZkCwUr0hmrwE4ImHV6bDI/
F/fTEZk+QBCTYlbMlkXhOKV/1CknLsPWG+GLs/1fdwG8rB4PRYLV+GAzYM0GSaE8rVvfE5/VJo3P
lU5AjwR6NwBYgIR/NmgjJVdEU+BIcGyElNWYXBYqJweUBzkMdce/2mSiWQZLz4CmuxiVE1dT9YSd
747ncgIbFexkrRAZobMFOveKZUFNsvZ6zvaipo91zNLV6xRpORbHRdw/JAkKke+sLLIIqIelDodL
LcNiqqqj8dU5C1qhZLl/xqhrD8j+tEyG3wo6vP7PLOZDkz8ac2/gI8b7/kuq+tfOJSnr6rMLcRW8
uC33lFQgoubuvzz4Ra6QLNObB4X7cj7N4Lq5h323I5AT42GKpaCBduHJ4eebmIUuWe8OMy+RxmBr
HfwH8MC9z1vDm2O7wX5FIrD4WtdupuJbBJlWtT3LKTm2S+5XdqQvTtFSt5Ijytw3cwV4gGh/Uy9h
Cu7WygBXRbxzN6GVYIO3IPoKGQKliz6K8pjY4cCqFoc+dItrqazKEGFH6HTjFpWmqWl/Fwe+3Zl5
XjrDhfQR2hVa4Q36ALoLbW1R0t4Rrx9eHSxZcmByuBJ8uXETxjDOdDgv+xHzvuifYxukEd84anJ2
s/g6ZVCDfqB9O9Mw6aByU4wySHXdiMvUpJzdJ1bU0NeRRBbXhzO2C0cATExp7H6T2uqWnrqnN3Cl
bJd6pLrbWTQhNB5fbIpGP1t7LvDWnZQ6PRH92xCBL7a3hMKnKsx8957cONWxyDNrawt9M1/HLboj
SaiGhfeKVuLceX80eoeebtT6Byiv0n5VQABkjgCIXnrzqvBtWLu9qUx3t50wcetbysjE7mvfM689
ca1EBFITpTroCLbtotR573C6DmeLj3aCpx7tVQqEUhPfm2ugkjd54dEv/tkNXQVsSBOr5QZhHliX
SGvCBwdrto3hbN/RUcxxTbXzFcpc4f6wbIuGf5GuCp7gbvQec1deZ9f9YV4phzhq3ag1KWlvXk4A
rRDKhjbBj8xt0bvkSfz7B5g/SIfPT0aRQAo7Yc9zFoft85nUS67//ZhWpM6HvdpP/+V1MJPKs0j1
OTwf+Ks8bMUulX33NG1uub1wk7fnl2git96aofbpNu22FYEU42C8XF+gnwWNvDS26ndmxYPXqoXa
P2Z1YIWUAvJi0uJ6aS1CQGKi9lakW9koL3Z6AZwNv2y0k6ov5pWB+a2VmgL7/OIp06yv06xpyB4f
0ul2/AoLSNBIkr7Lwh7tdp3HCVISPj6a7kY+4eWmwueyZS2URY3zHcqea9T1aHdY3BV86jq62Bnp
ynrv1wbltjan64pDc1xgIiWTKbDm7C7Lf94LczvtxSSbx9WK+/P0Ri0ccQgGpUP9JTncs5LzZDrz
ruNZxs5NVGSxenLc9IZNg7+BP2mQ6Gi1ZLwMHvDlMUEvmizGzvgxac07n6ZAXthwg2RrtIAPGfRE
azpiLzSXWWlAiCaYqyzYMwsuB1wo0F11a6EREL0hyliHXzczrFnlZtKS4h0cfqo/4HjRBy2od34Z
BRqKdwZbezx+HNmaNiEP/fbQMp+6nJjgXkgQKMBY/S9k6jUI+uW0yNlUnnmaIr2i3vVuujqWNLVG
HOai3PMiKPknHAfi4UCknF389GiCcWlEHwTMJJEldSaEGB4hOxKKhNT3elG0FVPsD7g2v1fc9FsI
Gjhe8RZ7qauVad5m1zN7llIKALgayl+eaSaViXT64Jca/FUfg0wtExiK0Y7473OIlB9e/06Uu5P0
/v0pfQCM4NOJophTsofr+AW2aWIewKbh3cO1m+Pk/HIq9giCN4dRfrTzYLIYoHu7YXESjZ6gHYsI
dMuoiptNTd7VihCg4ZM2QMObCWe6kVh3IR/hzCpplMMJvg4c7kxg6CYhL93F0ZW/yEIFDmHNvOST
/ePNV9mWCBq/TJa1+N8UzXisZK3rMyecYYKo8noCav5WsvTbTWaQ1nqGuv3dT0Qx0jq3nYlpEu+P
pHfcqgrbAlD9mDeywdxdOoNiHNytWY4Wnp10Xa/fAgUZZW+iZsMs9mfLeFPQClZZsF5osWbMCW5+
7jm8UPqdCRKoyWFQ4jxIk5mlYCiCCZ37QwOE1iguBdgCqKp8XPdS5dGgRb1egQwgQYQGiJz5sVyT
FZjAR6hkRIyUB6FMDSIHhe66lmQ47Vhq9t/A79WAQKiJ+4nKocnkIIVqOdSzOL9WveUi471VsoBa
bZJqNr/IAys6gSIggLSg8aHtONnRyZVpAfe1LXZ3+7XSd0RrII8r9Etj+ZbIm3WsmHryURJBneHK
1JP3Wph/VIUZs/XQpVr6WMawj2axOnjZL/npXKILsPSppuOw0mCgnVaAyxMJks9bZhA4LSy1IX9V
lzvwC29Uu95hUFpvkzZ5yx91JuovRms7+awqaojavmvgVjw8XFTrQDdaLwbIDPPaZKcLGYWWTdg7
7MhNOtzzygxFHWsNuMvhg3zMZiqtquHHrYoindJBH2FJvd5e3x4rmW0p51I2EUPfpvbmBQ4/6JWp
x7DmzszQgOC/pL2pRwn4RRGT1eYMAG6LlYwKeW97YsN3QBTNuO0bNbn64OtfL8rkbxCqC5EQOkuL
mWvCFJnFuW+HIDGrjiZyLdc8KlI1wlBfK5nfGaWspEGS+aJCendnjAkersn3htVKsDsNzjwXcBxn
tchTVIyV638CTuvNI5QdupM70QowSiCohUJWNLxxAKBA/KKL1xP9X8K0kVYuSW0kLTlEeVsSAc3d
XTlCJ6Iu7aN5HMgl7zscee93jhD6Rhuqe6Kov4TmG1BZKfUPVFJSSSYmDIKGEM1DhTIEfIbgWuZJ
dm69QrXTp7/ipDRqo4s8svz/G1qbvf3/vNUkGxIeQAhtggQUqAcacas474anVkgrFLD+k8kw92nA
HdVclz5SBM8IUWWzF5yvqMk1UiPbjBF3D+M9PnxbWEwt8MXS2y1k+zy+pZdrxYD+LOcLmDPKyum/
r0IELkahvOXS9nTqDJXCt/bzSegx1op5eUrS+Jqa7VovC+SDZURX2RRAWK9GTlK3XyyEadlMNw+W
sDBmPkyTnZ0iMqV7teIzx0Y4iTpM+t48gHXLUOn7+iXXPeMwHSbAytOA6Er3BZ4Svs6KO7QkoZT6
WlK1rZiSbCZL3G6mnsyiC5xtEbWhGj5z/r4TPtkt0bhG9YTIHi+iKyraTMpnUDoRgJ3qGm+iLMMW
2XoDmYWOLumKaVyp/+oB4YytQMv7iTbVKNbHOU8aiwXIaB+Qd/j+4RQ8BnJj35yjric5CxY7YrkE
SYEwvCYk5XYyK+XanpSTUYvRABOqL4VzCrOHJjOLBrJNb+AROgCThOQWFgaFgoCCFi0ufB5YYr5z
UyTWizExQB+2LHV7HyjhFiv4uVmSQu3ajKqIGSeuKs09KOiNYBgQtL5Z1u9iFrFlTrGAMLreII31
yLHdZoxQpqpsw920ok2bLxxxm5CGqTiIAnej65K+epXzzjUVPJvzMD1kOG16Hx5mOHHrjw9G8UND
94QC5qlpm4mq0qt2d+5nPscSh+66aj/YszFklz7N7Nt+m6hT+wo1maW+cHCtXcrq6VC9Z7Vhu8VO
s67annAicpDEhemEWksIBCH69dFMYj4ajYeuyeabgNaly3HX1g+kfYJe1CEUeVwBtZk6JY2cjoQH
mr6LM79trznunIiYpR3H+RJR1lA3pPfKpH2qq6kMQVtUaQiGjlubdoDBGWnL4/Fp4NuSMkobc5QN
37wDefL8GEFDluMAjFQqTnJ/Q3kaBy5G+Act2+vFvLb+SmprxzcrniE/SfOyfF4924v/XrvEqkR6
qbHmZijJdy0FItHoaYiYBT4nfNnGFi0V+04lJiyQDApcmevlKdm3wAzPi/FqpvAMqglnw00+xsOk
rivW2o9G9e5fzG/JmDwo9lCQd8AsZ3aIw7o40soyM9LPv6fLUBDypQcBvCH1BDvObmGt124lXdm9
G9OeXYK5LDuyyCoIC4+Aq3gFHBmG2qDR5kuZOVhlSe6SHTmhdm/9ubjuldFkZkNESGsW6644znoP
uCoSsDwH3trHHR9/Wr1moXs81IW8YBUpDj2vzipJzAmIA7S1JGQsDy4jqUEQGUNa/l+M3d/tjqvi
MYesey4OdzbCvu2oe1OVPyjLHpAQj6GxYudh9vcQFh33SHmE5RHfm8ElXIseotA1QVTlwIqjFN11
yGsjgKBq3RukLoUETqo9fyAZrlkUL5c8si9clyLy8gbxKsnBjEtwvhK1u/EE3bdNKNrt1sKB/uqj
cpylcW7Kf4K2O/eSyoyDn6Iz+Gb/6QfANRhvj7CuuYcYVsBnUOzkftTVr5em3142xhlAP4ACZzTu
Z6EOFOF2AKvkYzFCZqzD5AGuOiJtSrvJ6hAf6ZdHQJ7dPGEbJWTbI0Ihauj/j8Wri7OFvP0Z5zgC
Ql73l6CRatQnvr16wQonw+bup/tEKcZUFSSu9xztPOrFFaHXm82a2y3+vffMZa/A4oKOn/2qVkMW
MtDr9NF3LklcON+rjL3u8yzGUH2Xgs4FxeC03Mnjzj5QtND8Rvf8F+9zKFLGoGPTdYrJnIzoSLRW
gYr7YHygV3dqWOGEbXGlmMGmmaAiYiU0vXWZ2KzN/TUFgtT9Yr/o1Vdu+lz4pU4kaip8A93M6CT9
vtU5BKGK/x1KfA+PLYzehPIYp4Iue7nA6aBymXt9TrKaGbrT5AHnymIr37wjGzZzJaCOtlzkuzvH
1ZcnZdp4tq/pZHvHmo9Lna3+WWCBYtKI1EQW3xy8x8RY74RzHf7sPfLvn1ZW9nMeb76mN0M5l3T8
n3BJB/mG/37fj6J6NFE9cHqAtJCRw6F75SwN/l88YGM/1PtmfG1oHcLc5kniPZ5rWJIRDLeI+IMC
3H0kPMFsLn+DdaIIV9jP9WcvhEV3jULbQ6V+wR/OtlFITIRMX/vvYA+mj9nn8yHLcl+YcfflLf/U
clfEcCSooa6k+yVInEQfSWZHehorJBmpcDNVa5UnMBF1tnUIhkGZxb567f4aIiCIzDPtwte9EIuK
JylUxC4k4ndaRXU+0BdJ5pKnv3cPd2+t51rVn2/2LXPLnqHPrAi5im9CaLKoOH2EE+BwHzho7oPJ
i6naAQUavL1mAWCfXsIvCJw7nT4wWvS+kyA6QECyVM0uTi0PmfRoFdGngZNaV6O10PsoaySg3Zaa
YksiN7v7dE99zn8HjYyjreD6IHf70mRzGmaYdGashOplqyW0bSlPPCXP7JXybZ/M3HbMPtE94FX7
7EL3Qvk/btJwPU9kFz6o4RKDCO0iPeJL7YdvyqRCWMDOrJOTOIboK8pvPEaj6iyDoZHT7PxXuXrk
ezS3o6FQsNxOstAlsL7kQZqu1wSBExNxyA5EmIsu5uzPrcTKPodr+QDOumsrhj+K8AiyJ2vo2uVp
jKZ9mAfiEa+9zS6mpi2znzF+67o0gPch7nd8JyfSUctNP5S0VqHdc92J/ie+7XO309jnOFPMT0mE
+AG0nI6RB/getzx77O2VMxO1tcOk9oKliEgBXDaDCU4q5czw3FbaDI4uWlunBfJvt0hAWuuSxnWB
dOIf0zbtlPvXhoMDpVDGudQijWmFLT7ZwNRQupyiobtMwf0pHmZABL6fWgO8Yz2gRmzixcRYzb+g
G7COMG41QH4uOU7B6Zpeva3Cv4LePPj0at5Ev0db2ZisJllv8F/NNI+RC0FDNL6xWFg/qYloXvMM
QV/zdPdAWPpt4C4uABAf360iFBIgeAJZg4v1bEUnbW6FIpKVlwHaLX+Z0+ziZCOyg4mPcSeFcmRJ
IGlyExaDJC0U5GerSyxP4ZiWE4n9eadaoOCGL+S5LH/TEhI378udBy76HJO2Pf6CYFJA6+5WCsJO
rIPqDVLmrzzP6zSiJ8okyWAO/bMa417kH3Mb6XJEdm6XFqFZq/rFepFgafdKO274TS3NJAkb9nEg
weKyxNR1Qp03MyazcsEYI3Y8v2AxWZaI7Kwa8K33LtsMShnQ6GYhUCMmUf26oWdk1WfODbNOjkfD
jT/FsGQTjNAqQ6hPXEYHHsDK+08+lpBQ+YMNUJ5MLqf8MIRQGZsuN1f0ZKfNdMDFL9yzb5SfAMxw
UsLYQM2f2DcrrS7lFhLShGu9rbbuPQMzNhLPTPJg8EzFHU2+ZGxHsB1XSR/iVGO5F5wKNfQiWUIi
+T9Q92zkGFwCATrhNo9bNIu37yfubbpPIOFFeg+UeY7KCCl48fWdBntiz69SfEnLzAX+ATUCrUpI
Y+ZATdsC0Nj4lSU4J7QEirOFzJk3g+k5zSRvAwiS/zdLLxKLEoE6bPZe7e85dFLc2/1T4cHhj3ta
0VnFA0NCPD1g6O4uc0EjM0yQMNFebBeC+/l/p7x4Fq6WU8Wpi53o+tbrhUywxlbIh4U89IroxClv
FkiBNo/xQb7LcyjbGKfwBVjZi+LyS2uP6NoBDOLoPnWSHmSNdSXi7sTWDo1yvb8gAbTwMgBXruZ1
ILgiXGmliSIGFiZXbl1pBqZ3wwM+Kwy3szLuHH4EF1LLhbOznPDqxVNX7W5lv5bAk9IkhOROfMr4
KCHkVV5OC0dBmAqj1IDPf5IZXwKULXoP1YbqAardtLZP7/0Bv0AHde0lK8cSb9FCASWtmMwwN3kq
zYVo+odj6x34G7jU9xXunVr8IdNK+P7ZUzy157E5Uzm0PpGm43U9Rpk5e+bk6wUjcwtm73bxxanZ
OcbLAtSw6Ve2cR4GPnumgBUI793dYxLDN33fVarhKQEpGyWaTIRPY5bDrWvytEF9OL09ZYMaD5wE
pnNYcgYGL2psKyP4V7EvQjERoUznrqagNYv44K5Nkzd0IglmW3MFpwSPZXlfskQS62ShcqcGcFsZ
VUYGyleu0j0YnyamHJMNxLHKFrlWsCi0ZcKgpCwWONSKgTwHBVy6AP8W41mD+3bMt+ircMFHgVpj
We7hHrPgDEP/5/1Jmlk9/Pf5CugWyNPIQ+tD/2DGTCVZyUMlLaJZD9qfX4KqrM+L1c+bIBvFq829
H0Ww38Lhy+gY9JgsV27yoqftuazG9rQlzUzEc1ALRj+Tr6b9w7/sJmCxj+1u8kKOtNh+3tv0P5CW
J09djIL/ISOHhUjR6nVdUheo5eEqwBVopbh5qqVzemYPig9OcDM8kZje8wxgx3Q1PJI1sRN8fEru
j6rfenlnnLbJTo6InU39RJsfAC+rxlolfA8Ojew5hxACrahYn3Zmj9qyfiJh1pFeqesifk34Diyz
zGNMGdyStry/pyalBHh/z/X5hJC+VOnBMobOSVkdWWKAGraBv7yyd8CdCNO+btz7+Oj1IVSinCF3
yHtTsSFw5xohrK+w+jCg2zlngz+tSqON1fwbXaHpK0n7/kW8kQyeN8TEl0WiSxegz6fonLB6DtOD
bPESsPC8g7UAbfcqMjXGSvYZcJCRNJSstE6Z1AkjYlkDUeC0OUEJ84HnMbSLrMJb5aWsjBJsCMAM
v09xDFG7gkdEvkB77ZFfWYt7TYt+nzq5AgP4aF86GY6GZjR7wTkeyJd9HIAhcHLwiJY3cwkRwcGy
jNc9UOIolkeCtTEbJOQSYmzOF1cHlV1gOlRPjMentZ6MXl6WSpOGTShxWguanVlrzmxMztS4A2W8
wk5XP5qIkGxtKGh9HXPrHPj0Vez1f3twNiYKMZPXecYhxh+efdPrQiiuwBhks56gbtnKP77QdNcs
5L38i+oG0oMijMFqIiU6PFOOHz40iiqD2HR8ONhQ02XEONOAGc953JbQXbxNdt7RK92wG1IqhKEp
FlWZBByvZKPkgztzgB2osCZDLbqaK7T2+V81wd4wVI9l1mFUvawGcB42i65/ghI6URHsiD/FgnZB
fpCOEwCN3uHXtHwiQLyOUFqJmwXzCFwEFYwOw5ZkLzKzW8rEpCnU8iFbt91aUuCOblwqAUOSACWu
vO8VDro9hajhw20FX+aeRtaqDT8JpI9/8bGLrqGR10qwOUYBS22REdaj2WMVEp7hjzZP7RS8Cm8J
mQhz0Ptk2dfncbUiYXCrXaCAb1AmTyivnrvcMwfPekx42jYfRVsQ5QSRYe1IdjBsAo6uPihnwraf
k9bbtS0JvQdJezvb71SfkOFzsXS+XDV93/5KTo6k0se5wfl+TtDR2rqbUQCy37MGdfczJVn2H5fR
I6rMjix+gsmD1JrNDH3ZhbVhoPrBi3G/GHRmpuIOvJ0UCY/hcrUpobAwngjcAtBgrHs60s04MSo1
6N6Yl7AS5kAenOB0Kt7oiVg7xrpMQZ5ppHbjwmUuawNfvaUWQrimgCbauybDmnZyTIdkBIXZSV5c
9ecoq2qZUg8/xWVaPoPg/JC4fK+WE4gX80+zihUgoXd4bdDZmc8jK9LkhBpYW/J0AvqdGyFcwD/S
tYR3EQaTzMuyF/1A1kDzm4iLTSK38ovnVH0pR6NcoaDLnUe/XBMjnD8HIF+DFrpd5JHExIcdGf9W
95DnND8XesdDP2x9dPsW8dopg4r9CNfkqXEra3lL24QeOsAquDzrDEHJw0cikm/SKJq4diiD2Mfs
6yaK+MuUY2YGp2TzTO8eYQTt4xwvlhXjL5nB/c/TPTV9f4fA/LIbfd3eDqYXtM7Tjbe1SKD3xSm/
ka5yeVlhk4Xg/RA+1CW7+Kk/9ebAI4q7rV44qvk/gTvQpK67B6ugvXkee88CoZYabdvwhv19E2JH
5FYaZuuEND+JTCgbuK+32R5WqS9BMAh8KKYb8W3Zn2GPdLYoh2A75NAUQ5k6gwfjkHhX6KukImFC
YxBnmiIZVmHZGO/FlbWkZyIAuMjaKqD6zDi4R/Vk7fPcEEwJ0TGhHZ6DrVKp1OeBButuufn0c8ow
oGPbLgz0MOWwkFA+c1cf8Uyl3sIMwHCgvT+qhUKKgS4ssKLXSOubhRecfJxJ1og0vzRHVUU6JRVH
aUeQP/cVcBDgIcbCd+TqtnKU54jkvmG/0f/GmVlUEasF5+oXZwv7btrfWQHd10WwsrDGaZtaIPRl
+Uu+bbUaoR51yhSRhQuw2xNcB3MSAbQHUJ8oA6nrjBsLY8jowjpecJw498taQYWVvdP9n/Og7ETx
5ouYgFOv8AygQt8rfWHujzwJFJVgtZRQ5pQ7JDpfLhuL+T/2/QS7VflldZzWAVEjPMWZq720Lug7
n2rj+CboQ3Qo1uCngqxDfp+ixfQz+35mMft5+6QjHOBcJ4aCqHNRLeca0uVOmZ4I5McUsHH4vQYo
GMoqC81yxZKSkbC8oX5HIROVZmenbMthEI/pxmolXNf3EZL1TniRsKrQr5VWtSRdoprTaYlHaAlm
uPDqKfi3jMIFGJvGH28tie87V2KrYAaGmVpzoI8LGLH1THYfZtGtvRhBjbaD9s5A+HMU242v4hqm
gEUAJJAI9z55u9L/g+EBINDAJ2aTVHZ9d0h9TxacLwTw8kC+QSQ2kegqHmM81r3QBzuLOLsi05CW
mEKs+tCtVc/fCrvSUaAodSEcweHU8nXHUZQNGpI8HLB+r5yyjM61jyF4RGWsTF2th+POezXyp2Y8
SGJtkN/xFwJSUGwAFZnpQGGcmvPz0n9FMPB+Btq/rplkGoUaCtHYVhwUI/9YMod+R/Ib8Xi//NmJ
ypa6he6FVrA2bvSpeWQ3Pu3MUa4iDsOKeDQEHZRs8XntELXvCB6UO/BzacyfZ+rVR0GBclutJLAx
iUDXdOEaZJTKYDd0AoocoYM8EdVeYhWdyqXXVdWMMBDNL3sfNtqfBNh1Evx5NwWAqpaSSaJ5YTNc
51cOw3MpQrn0BWZrXwEcWQRrJJLC8xPA67ded4dHnNjzyqA9k/BqX94H0xz//DknjUOSUuHaauHA
nbl2fcT3A8exRpJXNU1w8bHUWytP9egWwkL93RMGK20xwyPArCGuXnpoQMREgyYk/lM/eVNYM+xp
0uMs5sL4dCD/r1CDOAVP6LpvWG5EiDx3211+j/j/71htD61cDzIk3MxdSDl3xxiX9Ax4tz/PkMJy
ESJpOC+Ghw9r5gvYJE8+smzjy6usOND68/yN7WM/pNg04qpdyCCxHmFnMnuc0ZqhNXImz2bcKarC
rvu7asTpd3v+NWWR1QAyUy/MGbMZIRONwoE+sF+5aWUoAPOqQrAMJ3yJsHgfIijZkrszi+kviuaJ
Mn3WWV2PDIGyG/Qif5dka7k1WN0xj8pZU7faZOYCGBjTZatcfqIQxTl6L2lojdwHqzLy2Ed4U1FU
VLkndwKkRcW1fkGESvkOTc9rHqOQlDi7R2Si2oAE9JYQ/WoaUH+Zhe4tU/T0+u+oQprU/n8aZl86
kk9AWcSeGA1xouA/wYzZFyzOx43Y4hnUFq/4JlhYQV3YSgSMml+SxRqYtG8YbmNkRVdO1ezKiRqn
qNYAHCYBmEfxs/YnBOODOrdvgCCFKpMh+BdFXc0SeAfPXldwd+Fyq987iMRMQZeys2FJU9jHwcFy
scshZyOXGvHmOH9/NtLDfqMglGH4kGYkELeafBs/g11mIu2BaBWpIMlshb7EVyo4Wlmewg+IqAi4
j27AT1CCPwSm+FNykAmXHTqo+RNeU1qrDKJtphYg+UuPr3DFC1tothM21nltfoJnv7+psjtvqmEk
QBcaJQpMnMEbCdTqWpEp1QHuJjwvVhlnKhZR1vFQpxq6C1Nogyd0Ra6VVg4A9SxBO01DzZY7qt0B
s6dWzahdnPYR3Y9iCJe/A5K+ih+QQko0Ar1hvgjDNDm9Jkb2KDz5DkVRh4kmNIls8ZFaxYRwj+eb
7tdSGVgEdM+ZWaEPVsllTfXGLQN1WWBEpW8jkewn+bd60oFQ76AQWB2lljOOLUNQwzQ0jXzhU3s+
aCEUHFWORM0U2U0XQxAf0pghjKEwbjH8HyNjIZ/H6utt43nzsfim/4Smc/BTMw4t+0CEYRUm5Bzn
H6CIgbGe7ZeEtdFJArJsyP6KjNGSExArOuY0kNI85iLd6rTI10igd0qcvHauDRX3AyY8spRW69+q
acQVLgduShTRkIPKWP9YC4Dz3Bd1YPydLIsdEFTxJ1vMKJk7rTwKlJOx9+0Z1UTScYEjWRJb04Wy
CycTQuLViBEZbTVj8sMUYYPI1YBnuO51tLGhvqPTLWPIHewSLTirOeGJ3CZ+6TJOZ7421GBzIz9t
xCLZKYuqe2x9JUwKrMlPzGewfkdDwdGFFEJacQ3hEnareLHM+l9feog15lQxawcTJMjcBRGcxng5
MvjonztXNRyO3ME9aklQJBhtuCDALIGdC3Rh/A4QVBnv6cRsOO2y57Z4kDQVA2Op2pdi01HKDTpT
kYwNzgaEtLDLfeiq3/+DfnypcusUMXPXtEofHwRxxAxuAlWEUv3f6a4dPVLZRX9LooYVDyeTnWAl
1yu6bJJ+nl9QW8hh4kU5L36A2FyR3CbudbJHCs5BGA9En7PE4JnJUy2tGIGaDLsYSwII4VxGclRu
09C/BNFN0LefMRW3/slyiAPeke+LOheivjvxxnVnBn76LPW++mzfCsao8H5rLgJQp10p70qFB0MK
XmUn96WUEZZj3rpBpAiIGs2GnxUwrSwEoYMdbfFHnvUopyXPFJMjeMSLKHFvZtppWPHNRj5ulEQJ
YRzus48q+RzwkgQGQBop8PW99w5GH16xmKKzTQWpr57sUqKM6l7nub4GxznHS7GiEQbH0cjcmtPk
MwXljdPoNNHnjRvCggDLDOXoV4kEDqVZa0sBDuNsZUAm3k/k/UHnbVruDR3Yf2iX2OeF32kplpdq
Q2IQMEYorbWpx2zciBaReKhvk60FYXhYlQ57C+tMlcdp1zaga5BLHWetwsY0gDhvIDPhGDpWbmbO
q3mKaMP8mDInGKTsdDtayMOLdmcN0xse2xnmiMyLQUZPNK4cnu85g2V95FTD/DxoWO++QyUkU6mF
7bFJRIVkipruRolV+VygGyYQcycdTyc8DMNAJOPaKYFh4vVqt2DR6X5jBYNxKR2CIvDT7/SRXY8y
rp8LWDyKOeFfJaakKM3yCBJkiBTcRLV8x9naRcISBcD1oPjqW8gmrpE+ytndt9svkU9vKmGl+rBU
4KIjW65LSqTELYDGqx099JNgktR8oPDclt25bmFU/xUq5MC7HxrVqcMEb0zNrgt9sZdY/HLhOkUz
kKNn1ddNymMhCVwYB/zrSbr0hoDASGBsrHvQo/mkWkfY8qpys2a1cD3SgNY1TkH2AYU0fkcdAC/z
gzS/vG3CA/+XBXhZu0TZxtns4kEE6enbqEXfJjv+EZQLQiqgUU4HN0m7zSdODkSMfoDLl0dypfy0
lkYMcJwfOibfGZAoYPo/z42+YoDYEFzzun/PxDrDX8kOqrxihH4FoubJiN7cp33ZmgYzsV0dzS/E
G50b0ZMKCQDTss3OWBs+2HhBpcPXjDYNgKBXOGGXsur8jsEYZoCm0/UxCEJpRTqfWX9LWM3msXRy
lApS94ugm56QHazI8mE+KC2yPZTtFL1U5ytzNFcXjvZSdr257VKeLvwmDPTpp42HIlSD9TXZFkCp
kR8OY941cbcKMf/44HM9a+QTCIXC1TfcQTDzk6+VIeUvYq2CMdlExu1RCbw2NzNWgSvOq2ffEBlf
dkQPYMOmVX96OHBouckdm8civvN+CXvrguJgmNdf43FscaMFicJIEOZHU+onuNDO5QDIGAhyrbx4
7ntD/HtSMOPwPZRBG28kvaSITAqrdcWA5anRQAtDeg0fKdmML1uUNLJ2yw/tvitQ+aEe807+GOWo
fMxWpSf6ZvedOuIy+58kImnO9ul/BKBfFDgrzqnOzR27U9U/DtJTTgMARPgdSI7iFPTCR8YJ7pFc
uN9XAd1K8GR/Opi5dgfOVhtDLlhFworrglm9gtRNPZAFWGicTbQ9Z9myIehyUuEOPj0kE2As3m/W
MS5GXxnh8Fqqb4FKdBJbpX2vAkH16geUqH7WDV8ya9ru19JB+jlJIkHLXHb1pvrYPVaEicekRQG/
F1NtJM2m9fhyQI+YiLgNKAJ2sArmXG7GbXQNddzkXFGdFSuINnkT/7NBSf2OSfHHyQHIYzXi9lwY
ZWiSjgmmk+f6dbgxKjCjLC1KZnqEdnU48ZL5MhQ+icM+iQAlZv/mV0ZfEFHmq5cCIaRo5Qb6B0FC
XbqiwXBs7R7Zu1kom2wJQtTeNsu3069ZC9WMOJ/+2PJ6XKpi4IkH54N5jVsVoTqNwQJhQw0DItn+
pP+Lu0NKmp/Itp/MdgkmiPXtCGaZycZ7EpH5Pl+3HW8X7VDSL8FIaA+So29XHuE4ct2dYR41F5Ji
do2WymWb4r0cN+V/yUvQs5CEpiqMa9QBhC/hsqRHwxyhlRDNRHi+QbXHLOB0Trx3Opg7AfpoYqCb
8KjkqPFsJlXsMfC4iYKAAm7e44OW8ikOI6Cb9Aek16UYDb6CZfQU3I4btQxVds8aSIrRQqUccsR5
4gVpzHCXhDgBarsWgtyfg3zpDTNmFPzTt+kppqZjAAFvi3n5QtyEXcb4jvOAJAPYsNlMD8555yPU
DCODSI3vK9VRNCKBbD2dgL29+B/ZtBSVvPZiNsWOERerrE1gd2CWAcDZSJCzv7OfzZZovMHCeLUi
F3ELCGcrW7Kd5NLZF1VQH7rHZIaG6ycUeyQ7Vehwp1tM+Bk3YKWUggrgN+rKdm0Ek7s05UlodaD+
Wkn8ZwnYhNLVycRp6alY+F5vPOKQX5FoLYNoG+z9CmQSXTArpjLIWSyO8XPE4oN1YaoZBx70H4hZ
S5P0JZ5iABkGOUSMTJEARtzD8FdntLwJ/+ZvdGmWDS+x7KFH6WH73xOCxEi20L1ZB9TBI/0PV/HH
oaWlOXjoZqHGK4yo1uCTefMQ+ZcQwfPmareDPTIm3NRsv9Tby7Uee7YqWYBzVqCnpEI5V52uj/Ya
16jnxB2/zt/3bLr3lp7L1oLO1aO1NC2WCXCJMygOLqoW7DXL8TwIDL2nMGgOKOLX7ndRZfLgaQnQ
YB35giY0/wriuf8A2TS22cAsPXDPwLpaoEqOvKEdiZVuPa2NoFvNkY2ktqi4Qdf4fipSRcjAJjzq
VVzJox/tf8DA/eZwFwcDkEjKM5lCU+skIct8cPxFRAyR+tdE3Gt0ZBARetu6FF9505VaDtxsvaB9
RBrPJSfgvu1Y+YI58HScdZCCnJMou4hSS8SGNvwdTpT7dFA1PjMvMpdZBcfqVDjIeajiLRVypV6z
BFBmz2+g1zfiGZK4TNpnJG9sao9FJC+gzPgmcwRAq9TWjO1xDkK8ZeU1tzxFUV4bLzKYcfOdKNGn
sVlZbG8UmR/XrOfkjhP7QhLn+cbTrIo95aPUnZkPi8yj8slmCgZl03hUNP1tferDZrICDRstnsi+
rK6vnyksiAM0kYdhePdyjG5KadI1NwT8JUsuWNy09tKTQGgqYwrsCeQ6h+PDRKR2WaHMKVHhd7D6
RFd+QTKP40rU8IHTdH0ebvH2fJUIDsZEp57loUjt3Kjx+JK9XnQ3l0+xr6sWT4UgYvxJQk363I51
/U2S9Y6jotzLpjU2j2R3pNaTF6xaJHQWOIoRcY/7aRZyMLXkpKPBVIVoW7q4eRCWUxfDxbDjnDGI
uKubyd+z4EZ7mCf5zAxEKxIovATFmHL9GeyPSFzrayGcA2FEdXjIiyMukRw7j+ZRCOkVVj7Jvkag
eMwUAnrTY0WSFbRrHJgY4/7utFGFIFIvUmghkhG4o1gN2aDmuDeFg4otrK8Mi20dtHnflV8yu+2e
+3duI+a+WQCgbfm//NErf3yVBfkrhfzL+CjmhmP6Y5XwVBksObSS0o7Vyv2tYt3nE8dSsF3CCLH3
ki+Xxhnz/M3vetEfN1/ATOhrIjfOgILd2wuNHzAujLciuDhXaC/3wAuDma6Y1wN8/fGFCVeEtx8x
Df+dk82hhPL0TWBxvHeDFx0BNIkaQpqj8rFgEExOVbeAt2fS+xStGn7llXc6FFKprUVYplu8cGFh
J3H7uojLVcmZgBxZmrO485zYTXPGOR+hepbTJRJWqJYWyXovGlbw0X4arMxFJAALjWlEK1DH7lwZ
Y1yQ+8gsrB3BE0zKBLw/b7IWGqIEk7V29GB57fcwyWC0Gl5AXtN+N/Jozkkc3cB5hFLn1j/LmZvh
0E0hgAUeK1j/Ch3dD59wnM8ZZFiLwyXkGgL+dElbuRazlitWilTbVDcggZzLZ9hihcj8Nnnh0ni2
/U7tO44Ql7AODD1FesPxBirFg6vshOjSnbF0IDCYLTWi8Erirbkm06H/9u2wY3JAndBLVY/dW+Y3
ZuEr5Rzqz5HQb9+fQqOIEM0vIaTeR1i9c65vwW0IfSc4fvteG75oRvK5QPl/GnkPi2pJXtQVkqhf
gnbHQ9g/qUCrNITMywPMLTZbU7S5WOe1APxNsWsfaYatYhkilhLlD36MiO4eLtjYmbEeRFGUOJ+w
J2TYyzcdUN4QjUXtSfSrkiyOwku9cUoh0c1uzVOO1cQ3tPe4vK7qSBZH0XSWgH2K6aE9MqHPLrbi
qAaCWhZgKu5QcQnNybCpN/niivBuC4RmrueCx3TTIJuphPgyHAY8NIhUV1CgmVoTqFOrgQm7/xrX
bIckz8+2QDWE2P9qsdgGKpKzyMV9griKBLy1w8We6UmGPzwOQqTVsx17H3blOHAqV8bO4zdNGI6J
V9q41WKFE4cB8By1+TMjiKtQvV+9Ggrn7ALBeW0ZXVAimxyCNSkAwzxsiXEtNbrQWFrkQbWx0Nsl
mQKU9RWsTIe1TB4Xz52MrKUZXDFW0Db4pYP/OJ23CoBbbdy+6SKnc7eThFLjZhHspQYiCCE6UH/3
BaYean7zwm8MvIE4ytEGAgxPLoBEg32ctwtYI5ed3A+3HJItdwqCQoccoxtRDKP6FBkpTn9gY1vo
hN53s7cuzAgBOubD+hUO2e/v6hwWA76nLBVX0BMn4OzGcK+oSEi9dMh6ddJFTAhtuCb80q2ucuFk
LCWIDThGujsrED6gfrGpa5rdqTZb8ExYskndHqT9cwkdu6xr1+/lZGwa+NKJqcFp8hmp9ihhUv6d
45jqbXUujIMoKbubSdmAKzCGX6Udl3VS1yMzFZ2IGtI28KeFKgOnQMAJtSlgT6L7dnS39b9LgVv4
Qpk2/ZCbS7U12LglWrbHZiCQw8Vd4qvXbE9zDCeYtBy2NL0Ckbv8o5jwu5oejZyVT01YTbfWO0Pv
bY3E5Qn1ZhQC238kcZ0pU/DDPOES5HWHz1jl3MOQDgeyWaEBagbvKS+sBrJCzrpOgL30gdly1Je1
CGhAVWRdrHqR0uyzpx5bZMW9O3tR4ooGiSpgYk2kQjmv19plywaQV9BVwyqvMT7l4Kv3EgSdwcXi
nBrFSWc9oP3UBQAtSrHiTiU/SgeUK8CxZx2ZTz1ZKJ7aAKZCKQFkyBN+CHYJunenPl+09wzjASsv
sxK5XoGOFkrxiqbOVcdlWddA0IEo0HYXYl+BYXgITS6+g83ws2h4RnJl3AEzj56bgd2sLNAqR2FE
esQHlX+ehnaggBppc1yU6a2SHfS9xBFsiM9nDp0eryoOTkgFvOa+VauGfEHFYiVQS9PdbyYneCFX
Pdp14pYlpS220i5Gr0E/t0YfyR6GRfqosLUGn7sF+jtjnM/8Q2UdwiqpXk4NFGd7NwTxn0o9aQ9O
Ok6xHZMlMthZe7vH2mwYnVw/GkBLZI7XHxpL2RIZW+GbpuD8mclYyEXPXuT8HHJhcoCoTlgiiL9o
qk3HBwPTHVO+QZEnxx8QDjiN/ytgU378aZQTHR+Xj3IzFjme8+ht8NiBL6QZaBLtmlnsH21ljY/G
b2j3ahZn/Y6UBnQja0mLBwUoSjXRKwsoC9sybnPdk8rUqnRVKO2fEWVEUwxBrsgy8AF/If4WPu6e
2TUmsiLfoOf3yBXdP2umsq8xuTPTjJeGPop/aOthjIkU/U1KeOUbdl0X2MWPyLAPZrE04FlowaVV
/JKETXh/D5/Ghnfn6u7QdU6CEgvz42CVKihU6ZOLp1h+fqqyc4GNtDsy0wWLIruvUilgFFwtCTP6
ILSp4WhyQ9uykI2NRj7jP3sztxXhoNpIPgo6u1x9ruSBy4EF6YKtEzXne09nRXTw5r9uBdlsorcZ
4BZvJgYLsrjqTls7RVchGky82BEsIt3Fp7MmyloAzf3TrRaWhc2a3mjmJHi2+wG+2qwCQGlrfyeF
wvKuSZjcJnqpqBwrHQRInAPzn5aUwgEijXP+zMavr/63JtVzZDJfX59OVf77z9aB7lI7G4BW7Avo
MiuemuMEWgKyvTugQGUtMgSRwlhiUx2n2QRw/Ge6vd3mbGYV02e+kAVT4yO8EMStzlK095CWtLCT
hQbkCCNwjhd3y3V1O7wckIUZvpY26bYkfhzVlR/atFGSvVX1V3QTinDwFZ+zXH1tvD3tx6z3srj1
HGMe3P3dYx03Y5ONsE6YkVki2yzF2dh4rnrzRz5aBktMo0dz926Ehfc1BdCWJhOLoAFF7Y5VZs1h
WAJh1+zfpZZz9PCio8Of0qyUtLvNvtP5biV1i9LcuVce7ddXHmcqz0IZs194FuXcXBfadulXpAbE
Z4fBopNuKsMc/UEocdq9+kpk5Xbur8wmaPUHP3kfpxlja/3vKp31ik320DPvVzjkukDvaw624bBX
1mHRYW9dnpQjhOJXQcsEB038/eICE5Zf8TKF68iJ36wIZN1m2o/IgQ9Mqh3GecJYZa3Q2qVYMaVw
G0Qgg4PmJgSr31ZyZ+4P2XQpeYpIiD3Mkf1+EN7kd70dBXERRldkC//SO7ugj3u9Y6Y78w/qPE7g
QOEk5cQAUrG8r6Y5N2gGJBLL7JA2pDJ7HwZtO3C0Nnzf+i/8lwMbkgYXXzM0FUAMNSxirw3apNS0
7nXik9Qn7MOeonlI34HQ6szPlijmTS+XL4RjS84RVSjTNE3j5q/zQpKxVg1bbsOXaZwXkUYICuHu
YmzJw+Dm11QxjVUA2XoooELCMqKdNhtOfvPkXMN9/iRKX/0BuqCe1upjUNhB7m9wTOg0Bjv2KkTv
/BzmCMbfrPassv7R+hUlWexbKTPgFm7TLv1CbYDojaHJyI8IkA0wf/Yw+EQkbmhne95ZG9LYG4iv
NcPTv92cZ0Uyc7mkOfzZSRzeYHvKbcfQQuo5k/lJp9ubQ+gvoSdz3ChJ+hsP13zcmp8x7J6yO45H
ysDpohnFzaUH0SgXokBEd8hyrEWT1YNNwbbea/K1Yqqm+Z8Htb3AewST/XTdA1AErpf8JzsX2Csx
z8oc3ht4FeGspgcI2ztLrNB46KePDPMARwpP3Gmpf7uifgLIFRIBTLjQqYWP5+6oFmOw+2KGnecZ
HDhLwMqYY7FuUWRyAPqvaNF+2nUoag6ozVUCmrO08DXH1LEP108kRVOYhvewHc4s78lm7x4x6eWn
brBeW4pbbBkV+CCCyT5ep6MRi5PYD/xlSZAmDZcIX89Ex0LdUN9UxrDq1pT7dif6mij/fOtg4K9t
EQ96/HKOcmC3rVu9NrdjkvfDy+6GVXAAls7wMIFPAZOzpYXZ+ZDtxw52HTfeqAlVtSbC7Dh9sUgg
eh9EkWNfmaC451MS1ebvlbhQk4SGVoF+2p6UJvJfmqeYHHGmL2cYy/8Cs0vntgn+1nK49RgfdVj6
9p2kYmt8fzTl8aTzk97zBamOs2xtRqwTh7sHrR8ooIs1DHnYIc0hmpEw6FXIVPmUFRRFo7Oo5ocQ
Q+rCmF9BE6XjEBYFgzy66Hoc3xbDNAGWA0kuCS3kbtYveDquk/jY23zX3zquHMhf21A38qf+J1Ru
OI7PtzWOK/wTvyJBOOTwstz5jNTb+ZQX++9VJ1k9PauakDydjAJsTVRq6muOJpY857AaOTCP0EMu
++dk7Mj06Ev9FUu6cG0mh3vOkrqmKtryPdRhRvKj+H+ZN6MCsQ8tm6IjUe4Sh2EEqBy3ja4ZJXh3
UYWm2YNW0L0vI74tOgyGI6g6RAa+XZMQHtf93eQwj7G9PEYvOEvWwLm/PHwgt8Js9VNApG5mJ/lB
TCV2hbHA/g2RO3duvxY2t66w1R47eHifORJGbgEmcjDN1GHx4cWgGWwITzBSxPi76vugkUmK8cMU
4ALRQ3uGt+4OcSJyy1e0JM8bN5GrsUZ486JL8s4Nsji81K8a50MhqmhZNEifSw3ohGk0OvFOZRrj
3JlyYjl9bGaPoX7hvjEpBdquonxY2uLeCxm8e4vrIBQAdiJD3IUdYAidEzBcEHQ9kmrMF8v9OrZ1
oJW4if18dO3XRqcuvlQx8kaelCJBh4qJ2LyNaKQUBSR7bjSdPgzfo92ee5eFJUqonUlaGIfUvI+w
ryDHRJQwNP0+N2Nj5dU0kj7eiHV2dqShFfHMfmYc4+nPM9qxrwH7Uvd0kOLuMlNca5d5C/rGkmon
sSbNzbRXYI5EgnCko6MWDDl5yudTlOfnovZ0zoYy0vkUQi9jGQm3WVJxNmLOR/iW16/cBbkp8qzj
XqQYGk+xxJeNQXxFnLgPjoG5QTzumLbEZSsVx686MDDVvVI1cqIF3Csu9Y6Y9nOGg3R9l8Kpbdi4
0q6BXNSfCdmxCxXHLgHmvTwF2n7kuCyU6oOtHZ5HoZIYa5HqVZS5A5LNFYWjV3QxHWQMbF71j2la
znvaKpcHppXp4ys6Err0tv+pI8thlzWOgj8p0Pkjo9igJK6kC4le7dktzlglEnJnPziQJqWUekLi
MW+Te/9gRQkESHNSmp0YO9d3rA7NaHHkoek0E+zW0y0EUGMc6I2Sr/h0G2pZcxprEQojERjwC0pr
HXWrmDubZkK+7BtPU46zEBWss/tLvxF22Gj6J2rYTsL1I//7ZN3ksaMG/ACVxI6BY9MVyWp8sWnb
eH+IsQB1FCjOsCqdYyZQo0OdBnGKQ4+YELo9IG/5OUR1VWyOhj6vSkn14l5KTezc5y/wmm+/dlz1
zJiNISx46bHQ5tSmSve8tcF7VdTaxZO1bzjrFwinGCe3Y4Emzy79awPEUVs+i8YryAZfPma4XomL
5bwgMOpbCps28G5LX3GxVr6qMwW8VJJxGesZG2w8QAqrz1lNegw9mLHti3/ZR8XWfgFB4n+YMjUI
LhD3kYhv2bDYLjsfXEEMRkkirfh3IngwZ5Xdc2urRVCypuHMQi8VjfoKb0QDVXVRV5fG983P5I1a
GzJ1aw3bhb4mfCBAIQNCX71ROk0Jiax8dMk3FjUPhgWd2aoAuwSmfS41aBwBVuQtLS/AOCfTcCkl
AoX8qNZpqeaR1HG9UEGNK6Ja33MU9pOwZSZwnCUb3XTtJb6oDO2l6qg/jMNKvy7GctGHBxDPPMp5
3y4ojV1AyxKSOa0py00d74W9GJVyi+lrKezFNuh/LYRLZ2qifbFAEnIQHYuRYvJ4F9V0ZYI7FohT
5bdOaOZxvcNSyZftF4u5A2dvaGI/DXujEIqOR55JjFzg/BeyXT5thM3uI8KNE3LxiTMDxq/EHda+
dZUiQX46gVpqJG9lfe+HVizhg/PVQrzYCV6iOxbN7kjxeWnf3V+4LH8d0j60HzF5wAIZNLuzEXYy
yO+cYWhB5Vk+CUgt6dxw+tJ3+fTL4bN6bNLSEl03v2zC9KORDkxf5mHsWGo0JXosafDGibQw9PEH
UqcVrcpUobwMRFcPxqLNbdyzZyZ1EHwdYNY4H2mRZiFMesIwFSyIfA32Ja4qEUVstW0FwwRr6Qu1
xsdkHiVpGW9YbJwPJugqvn0JzqXVnAFZyoig6cagbgLnGqmbt/Sdfnr+C6k+NMsC6dmZXAmc5ZA9
LLwVO60Ln0tU962vOHvpXnMHlQ+HvsxUKgiMJizVt0/8Pxj+HS9M+O2n6WfOkrPNPO0r8eoEZatO
DlnucYZ9dBRhO9vCXTBlviU0z1Nz7tz24NcpDAICV6BMBO4q0j4oduEGNrV01Snh8o4ijSWKgUYC
lwfiI5WTCriKm2oTp6bOHocqGfitL60ZqtGlIm3NkHJXD+VRvdzNOBLTE2ip+y9+VrI6uqoa2kp+
jx6JXmg/P2iNV+i/QqkQiTQvi68oYBfftlV2YUCDISoRBxikJXUKPrVacSAC+UNDI3uBVSSxbmoN
MNf6xFhc+mGDTHPUJBfkOZSlYO1rru2u404qfdWbzIztlyrMfD/stHYFnSu9DzzquuVnJyq+5qKj
WmxlF0QE3luIcZ5bX7dLg8H6khEVlAqX0Acr8TV2+2hyLbmlSic5DbGdrN3lnYmMuuxaBj62DK7t
tvN3lwm+IKrdP9SmgnS0hkO7bCk6gSH4YBaNxjGsh2SmOscUJukbu/NEYuCH27uD81JCqvORr7X9
KDrSJUfolAQQzq5OlTC1utQ9A8n3QX5ApiOKby4hyd9fSuPIVGhA/kM63/l6jKRMs6fNK6tS4/tw
j1FAQbH0KXBVcq5iqP0d42dTkhczsJW3yASeMv05U/ZmCtglQrqb9h9tZtCPGJXqZj0ctbSqdzJf
JmicHUZHw3tMc3fp3hzKoI3vpLWG2tkwt7iJOyUxrls5pq7kWM0+k5ex25PADrwjkVxuErPcn6rJ
Dd315Ivd4TXua/XhFehnLVwKp+zhcqspmRHIXR56A8uZQkjIOtfmvYJ0IbrlwSaXpEWqtXVk8Egu
6my32D99eN9OukYfRx1qgyI0LJ4grSfW3NCbxIVo7FsiigBefm/YdYGwr+EKjvuwMZ0/yYDKGCyT
DGmX4ItyxlPk+q+VTHqUP5zhGiHHfVcEzAuyQ3Nx03gDwO+wGinZyykpwalD9EH/dEaCVys4IxrR
XRkKJ6lUMezW+PnXgRNcLO4EzPrlRW/MuYBQqLu+k37F36ZSDydmzUvb1VCMm3HL1ccRJNk2Jpz2
ufBLzFYq+XuFflyIo7OsrVSOnh2IcrFpIurmXoB94WGHxb3loHJrYawUG/g3AEzPO8JFjQVEiliu
7PB4bumzqC6VTjPjMhocWyw9Pg8u6SI/d6qSlUFcGimKzR99oMbZUCfnXfOUUGc7RTNE6syqnSJg
tcbOswndThtjqsES5BekhUx97mwHJoKq1STKDuMg2Vhn8HXR37WLTFVjVSjVsRzK/rTkRzFrs9hE
EJYddVx8XaTkQH/FsRMutGM4zGV8hf1Jc1es9mhYS9mWF9LwW2zjyeSyk1tjKnJm/WgsSzMPpcX+
qJKSOTbGfThfAZWEvkg33nFPwvWJRsNk96FO4VN/chISA+btJhvr9twzh0Sn2yz7tw77Ve5bH/PY
3/lDJy6/I3dwOhiFsWxm8lQOb+d5HfxM//8DT5R8SA56aXjBvc1IW7VRc11RrtqhdnJGmA6nDpSG
9Y2wVTIHm4fGWvv4gWMbqVEJp10KES0TA2MU4Lwd4YztXiIKznmNHhjIAk6XoGuhODkwN19+3+oZ
IC+/hFgygijBcAgeThnkWII3fR1gEDVrvggYbWCh0dYsDOunxyspz8jBMVb6naB2J9V6iO/sdr1s
9o9h/d8cmUeAJDBl7DAxxFbImg+vwNOgMxaflfp6pIjazwOdpCVE0keMsAzo8Y2qCNqE+bF5E17N
SvVk2Cnv5N6vbPIEUsgSMReQIooePpnqaS2Zmkp/GJ0KtCpYfZhbPuH0sa5ii2WdEGxIkepWaIXx
DSRjulptYh0wgieSCSBX7bXARYuMkS82kYHkCHSFT9sQcHhI732cT44nD1Khs7NcIjGIrwMwVXUy
q1oizK/mA1Oj0mRywCA1EIkvzPXs6DeP4M1b9c3nCEkInxsKN9jZ0vnfEY76EulphZKLWJx7mYD4
mgSUDcX7P3W9BiHaoro7ItsXCF2A/xTWY8q2hQkKHNMfu/+FTDSKZYpnRTPYhZcmLo4wn3HI7M0H
EQ1Qs4GW+x/6ZDC8whihquUx+PKPg8tk71CCwnoohxSLBfuV3p0fYkOb7RsmtsVhDTN4/MpqHXy/
PO8P/v4JYv4MkW24j0pieK1UoeSykkwdJKdK6m6XZHZ8Lz1ucokF1iDwRRQX9GX163vipjS/Y+hn
zKSH08vtWpND4Qb621E5D17N+UWghWcMQYJolI0fnxnnwu7413p3gR1aBXKw0mGGAVEBOQEdLKTe
taKLZkluVU/iAen1SxO7G6xyGhymiyT9KX/sfoTROeqOeJNmShQ+Q+TMJNYdQqtS0ex3MqDCQ/4F
+SDcEJq6RVE67sQKy94uTPpqnSJdzRWPWlpIo8Bbbguut891LCuJajc3z4vYzDDSOtCHxIGivQIC
2GmjxsCs9i97Z3sdEWy3nUrqZMlqbPeyzt1rFYc1IZNV2QXyvaJMHHpr8em9W2shQfKgt1GxDjO6
gC3/KRl25nyStUAtEGlR3dzSWp1Bc/zKA4OIUJO8dLoASKKNNjxAdEsHdO5JHWwaIPWEoyqX9ti9
L1sBZ28nx9smLHNU1zKXjOKli6pyuZ33dT6HowTVe1NtXYZLd/pkrDBl/kRs0xPkkHWAJY76cyYM
9OItWnhda7UJSM/zVcrjqUHGuqmmsAcfB46kDf1HtESSF1rGbMHJ2nBQkZ+dkTtabOD3CHS1Pg29
FLRpGG6CtGYE5uxaObkxHAdL/Zazv0tnOEp6h4nRPChs/Br68TqBGIypq8IccLPqH/+IMRgSfS9v
70uu5GDEu4d9TWqM7Gpzdf1kBucWDIjSxC1CKb/FqkAzB0Vl50aCdkwSEc3dy+U9D5d74APYgvQf
qRqzFZ3HQdlDxfWGe/m+pJKHV2c7bVKUQmckMWmEBgkO2JxPyGBVDKcMS3BFmb6rUdKR7YKtbI/f
kN8BCoyAK7FKtIHdQ3NDPKi5ySm19J31tgGQHwRIBqUbQEUs0H+1qCa8G7gePB/z6exOP1iZVL5m
06rhqFOopVNlATycEO/sEzssVg93NlkhfG5G0VS3ntGOWnNXfFtkT4T3LM3fmnB7O5CF0Avk7qoX
vfoCU8WWXGfOZucH7ByQ8/AzFxIVr5EAidlwmqkBhCySSqWA6ToJs8b5J6aRYv/x2zJx8BwA8G4j
fLSkRyAPiuuEvvr4xOx634TWdZIPCvniCR8zuTZrGP6JGT8iFNJz+wVJtiYLgtLiOXKK4ygZr9XD
ZU7VMns7Clo5g/b87XdeNW/BZZ1o3Uz8COVGlUb5iUDoPWuEkveoHcfbiopR6q+amrBGs3PraSbh
0bglVvt90SZFZaOTvn7g0E2Vf/sJwyKdVcKynDFGc6rz0G22G3jkM1TqSVs3pq3PySdGBWO/WiVZ
mM3eRD3UPtcHI6HLeabiuzrGV0P2lqXsLACng13VrQe1u/LL7NNBYFjWc1YZ3v4Ng8PBiPLd8Pwz
P8IT6z1v7nJOYYcc8+l2kZjdHvf2uiIT6tslrp6+g3VlN8IgB9dLzRWD7b9Qjss+Tgdq+v1ELscS
2150WaWxrbZiZJLgqm4fL6G4K/YilIFNzTxAIEwUIrl8LcKwamq5PBdw88qcrhxvJ7HKDKvi7Jg2
TR+iq0J6U0plCzvifHQFhYrct23sP/W0uLMfDAgDT0E9lwEoRAlPjQos2p5FVyv7QA5+Pp1U4x+f
hwGED7PCeNp8QCuPd0KKHQYKX2UeCkdW5epJxs75GvRlFWARRU0YJXr5cpa75Hp0igU1AwK483s0
NtaFpssUSnf4/lmByhkp67uuHejp6AXUPdgvZmeRCKPu0H1WDhyMYrkuajM3IV4M9fPtX1YxqDrL
s+JVFjc93rWZ2NT7L1O1JzvIZpMsvlLvspaUgSGrAwhMZX/bVX0fKOlPoomNaaeUOll0rhpF2Yj8
lyCJYEJpYlnAaTuhXWKKh4tL3lcUF06JqNo5scoVakbJECD6Uvh3//S9/FUJKfJggxd+8JlKzo90
v7v6nzPUCGkO1l0z6P/rBXWsLD+BCyxhZnKDyuY3ceX6hG7zqXcQ3LeOP9iToHFor18Agy177NLY
ZoDoqvnON3eIue2ELCl7AEGOru0asdTNH8Fqy0RRD1iR9FghWRODZsvNPQdkro0nEuzMxcwf4s4P
WMbVzv/c2dcLsWRUzuFtEKxfUorPjpvL2xzCR0J0v9pZ8rlDCNCR4sBNtylRX/JStcfMraaXJznK
IRRgMoPfWus+G0LYWx1QcGtrVOkS5fzkL2euxP8ObxMTSA5Umt6EfN1dIzlUo5WzkYWj6PrTz6Hg
EADk/pXEQxEKe0b3WKGLOsIJAzY1f87qqsjwJQdS5IK1B+SYByqDmB/keQvjdvLNQjv998f0TcSY
8/DvIbjBWDZquUB0b3RfgLmWRGeU690fw5ANqpXOWoeGW+eI+bnuW/D/d2LtYUeFMwCc+A/YyoiE
rqKV3HSYJlt4uegzookOuucY09b9MQt3rdAVzM5LBiEPSEXY2aXWSCZj3HKoWNSAT8WZIo8SUmpS
HrlsG+cueAlC80E0OuooH9WeMjVvRhPTq2wXRbeJJsQekLgPXBNfweuVl2GINe2XqKU5dtQXkld3
4SBfSul0KXffvr7tsc6SNAGwj8nzMlzn4Ud1aW8uzCz965vNmHlCAd3mwbMZFGQHZp+47WSBLMe7
3iK38IxjDqde+RLlnpsW4dju/VjAzl9eqQEiMNIo4ubZ9xNm8RG63hxvpdzzDuQqb5kZwgb0KcdZ
uH17RcIfuRIpJIXQYu/YgFbMlPMl336c4DNCkH5pRYMB2dWRXQRZ4BQSRHiXnj8k4MIPQCx2H9mI
4c3XasMsthFlab1OojT9mh9Hox2qZ2zpCATJH8HiTo3nVakEEwg3QKBmgYf0t+Y7bq/sZzMhETsR
WuLmiQeY9n1hRX+0TlItzpu7eUrv/7COrGcoY+gbeccHj0HD2Kc7IOGo5qlVkQV2BCqPso5itxHJ
znR3oMKng2tttYCZwdfsQ+QlyM/uvmxLk3ZL+JDNRZDCoWtGZupGlwcAVaL8yNRdMkCmg7VM10xE
fGEdlSPcp0X1sPNLGDwmmUpNGLFJTRJzDfDnTzdQyxaquNNpe0U4Y8g43XTKFV9IZ9ZwE5pXtX39
sEav/eo/cfEKFzvowktXnZgBwZ5VNr7ensH5jslwjjrdZP0vY4wS2YKgu5LZ9QZHmHzavHPLiou3
u0K8fKklGtNjxmY/zjLOgFEHNMolJBwblvEDNVVSL5sb45rRyPut64RKwiIDXlV+sgy/Q414VXIb
32z+wKEyLNp8nkGBRUDrtgtgsPPrYdJHGHRW/lZCyN20DyfmzJ8OP9CQ0Tto9lL+OBoh4akzkr7v
pwagegeAYzty5y1rPIm02YBvyMDbX8mbueK9Wo/TTvs00GlrfO0fFIqa2kBzGqu/17wmKqFKrPzy
tgPZPYWQ4ffi4yAEQt4Y1dPl5PG8jW11pPxCu4LJd2HdIXPHuZXpMw1yEh3jKW+1p7R1HCelt9u6
kIpG96bv6vewZJ7wiqhe4kVIjM2jljGBvKch1LRD0JNSZUvdxPnZa4TzwC06kwWfW+J6OOMHnytg
kwgZSpST3zK3fRJZs+d3s2SRxtKSm/4v3raoKmF0XJRfmKMc3em3JSeJ9wwE7t/VbhRA53A/ySL4
b/Hs6Used7n/aebv2Yohc+WGWnfjf8P6ZEgbyH+N2ajONrv8noEPWW4rbAQPiS+adMTIWgFAhxs5
G4tyHWoJOmp4gAaCztvVWu6J9HM1Tjp0yCJUUS1wAntFazi7KIVMLj4gb0JoszBKeCayaL++ikH/
ygl/rSEVGekV4bvBHi+PfQDIDI8qwwaEy4XSaRT5J3ooVStMcAUe8R5NzdZNMxYsYITQz7s3DXTr
FpkVLAaNPYZn1P0CDGpvKi/WiQdYCfUfYd65ex6/VK1hNidba2UgxZk7D0r7s9IacNtg5+PVtaHH
TXa6zZgjFEa7cwVVDIvNyE6DrEJO/7QNEEBaTyVAoNOyL6GTYkG/kU0IoZRgGMAiPMdGCRXGIkWc
9oWs2dvkDGc5/6fqDxDJbW/jt5IEF0tXx7Zk/B/z9Y7Df/Y4ocjA4cbvw+D4lEDMOSroKFHJ9aPo
xChzCCKNNv/v7LFv5ok2XWlhhlIe7UzUuDUg1T+6jBmbRGKdQWlOvGKgpZdZExO7RIAXKzmSa0Jc
eSOQYHPk8zu8B7D/FKwFXkxr+foyyPIFWOE1fU2UikAoCUvqPlvOTzAi6jzTP6wI6FiKWVo06N/m
CRQkwn+LN67OjVBz0YvTx2MZD5LT1XZx35ftsVsoKGm7rfHX3s4ocJrBxIKvmplq9EADbVqIe7Ca
CF4PA65LsY0wrqouHrQT8bBifBIW496Z4rKkDnSY3Ysj4jq9iBK6knIVAdamdG54N6lyNfAifaBE
uabEuDUGvzpZujh4dB+B4DLVLBelTIAN4rJ6HTt9jxUQ+JsCoZFfdecpa3NxIPBU8gyvLbafwCjC
MzlkUihjvis2oIyqu9fFDseZ+n9oDATdfHWlJwu3VyRkbikoEeMLSaALrQjPefv4sPujoUcspgUv
WCigCfVJXI9TJI3OM6gVxGAtuT+qWa38feOe7Udm5rMLZMDujcNmm16Rro7ui5R4fR1Jl6yvBXM9
T5fg/Ha+VJ4HvtlmbhgcfBopX4QiKgBy0+NEUuiI2tn3RNizlG+FgLRqGkLEsy5G2HxnKPDMdqhS
oCCf+a/Pcpo4ewIXXzasp6180U2b5rjooXjWMoSLLfOAspKwUtCV7UpgqekYpcga/g+8JfGYeHuN
uXxPN5aeUlLOvrOKVIcqAO9ZzR7nydwFIqQQ0rk20hS4DY1hAQtFGPSG6XrB/AMQZ5sLK/Uh5n1c
eBUXYbPFMvKI/D3/kZaBtAqGeay3SIwnfP0zflpNGFwYcFMca7TkMZJIVaPhhYVS+wI4lQIN5BVq
m3fD/8ZM0VoinbLKXYwJ0z5Rj9m7agRp+kmyEIrh0rGgD1VPKO8lYn2KQ+gZT80mP1DZQq+vCzwe
gKMzaaTTUPYpvje8i9vN/WHz/A5cBayhqZXLfXofZp9IEuCEHJIrIQzCKMCZijarjArIFtw3eI4B
oyKmG/A6+5WyjSIzjLC64vrtk5nd7vtdkcCs6y0qSgyBuyJqundSEfk2+jUzEuHonvUBDODPCpNw
B+081PGnb2leanY8eX3J5hNK+aJZ/RHCLzrqxrdvN9LpWZQyYv2XElU0Wfu9U5/RKCybqFwrIP75
RCDAgJOZFG7qhSOXKwrJhh8IUOeRxgRxiJ7Ti/GAYQN7rOunAYBYQVyZazhQdYyG6W6e59sf9Jsd
A5oQQnBKmeJyUEeKtpob/KVC9FyavEvf6rXiH0D/ULtQx6AcDC+aBLnul/57V+TUHVCC+WLHheuc
8gYQsbDXCKJwHpB64ynLuVhSS5POXuWwH/591Wv/C/4k0M88+9I9OUPm2LTxg61V/KGppEzrCI8U
mGjppO30AU5666/txbOXTsDQ2KgjL00tMtEewu/DCbPssobnwU66Z+PZyGZ5XYX8nuOu5v728xfq
rEsfIYKTeZkpUZeafGPpgXyWPeq/FNDunpjQINCLF6X5nP+vb1C0fbPq4eLKaeIMIF0Xnl3YcfR0
1BGgsyeeVcIS/RKc7h8FvBg4+MKUfWvlg854NSei24UT6pTy8Jh8SULpuqrAU9WJQxKobnvLSAIm
BtfhURFRRB/cQyJBTOuMg0puSVNMpMfNeO/TH15lTFptmllj9hhlPBNEm/+ihNMzPPLGQ6RnuXkJ
dzBHptLVSbEwORYo8Fw8OHRH3Pa+/3ZU4lSUFzyMoU8kSwpKGvGsEG1aV3J/uw+/cy2n+zPESc3D
wylUL8FoGLBXfMPCJ3gKIwzo86FITnbSjaXGl7x6FEF7FXvSfYlvH8jiFQDQuwBKumpsvZiWAv3N
Mt/x0HqMDm/looy+wUmLaU70eDvxN7W5oOlKgJJDqPieePlGvy3Wx+x9qvO7OROl4PbtbjV+ZhGe
A2DuYW9Zi7psrPeOTMSH3evbDcP0qwiiYosQvnyy1VtJ7InIN64FUlUScuU5fYBdo7AQKJkw3nuA
MrAak0UnemXwhb1tF2BpWc5Va/ki2ylq35AiaIWEgXLA6cDWOyyMJODId9YbQWXamhuAo7y5gWIA
qTS5SedZTwRSZD4oCIaaWWTTaiTYStFyObqZlb/DLDzZYKMaE/b2BvIZYAMMxPkldWLhwfaWiPXs
/Xlxz1yvZY8Uy6dagj3pjyRAsl52zkrDoLFrpRPzhp+AdtTpdRZsezQMV3so8zJMkVNyZYPuu2Ki
EmnzbVaAt8q+oRdFY9x1o/CcVkq+3XA0cRCwBEhEVTafvsPplnBMuO9o0p19lPU+0Koq/WFOv5it
Rgpjgv3w6B+6kNj7lvLYRpk+WIQaYwFSCSKRa+YEsKznW+mk4QifyhMhhfuhdbLK8kBcxOCjqZFt
5BvXDwiTPnvRQh66f4ks71y9Be8nz+O3f4I/BZFhb3Cc/GRxkhSvvVxSt9bHxxgefKgF5K9sfxMs
gxWMCX8LsUdMNjagJ4xqJzWuI+NhLqzehxAYxVPYTrQ/T2F4k+pkY9Z4EiAPf47Qk7FHWB5uAjT3
FWNj7DyVNNDiVo/RbgCxsfURnuCOHYFc5chPR/OWBdwWaK6wavIFVg/EYjuwf6GoLChj5RotOZmK
VayyglGPAoEqupFTToWG7TZ5b+MZ0mnFnS9PJNGEHsHrG3j7P7amhgOg5RQZijv/xUjvQFe4voRF
xedaFhl8cU4LjKxs0QKCVFpIh9Si8pfKX+p/uguEJ3DHz98Zz/twMjDlHuN64KtnNM/InuV1814T
DTQjVTO3211TA4CZPvMqGVeyQYg0pZyLBR4yuWhaZBn8/HolXDvzUkDmpuf13cHxDFcdQ7256gpm
qlvmMp9tf+rBXbTl5w32fpD43EVsMSwN3zdPCDy+qPtRX3ziPV9MuwAROgdYuSWxrHz7kY4UABjS
A+qx2s/0wt/Jfcufim8uj1Qz+/PWI9M0wHZrIWReVbeUPuZXn4gJo1NGPECJPkJ74D2S6kkfromI
W5D/KPFwBBQUqg095DXUqGM5vuiLTPMVQZNMBCb28Pj8UBREAuFGTUUvOo+QSqWBQysdP4u6sfOy
mfKVOVWrSHZEGvbWYhJIIt/TsfpVBohny4vlsSGpAh8US8A8yaR4DH5LJ8zlABdKZCZuokc+1BAT
9EUhEHT3x/LD83Zr6RXedisEk5GLIBfPEZJJUHjRJeih+y27xwSMT1RUKJJeXxPnrgOPIDI5DqKz
jTv3SebYY5P8SwKzrnXTFNX6bKNiW7IsrXXcY+rkzMz5u5DneMn9Z/pHHV7QOrnVfsddsAZThMzU
zH2yir+vKsafZXKVjwJuJjVrC0Dp8FTXrxjAhDS+e12t3TzHvnQXFypuLf/XuactQXVV2A34za4G
BGJ+8s/ZMXJ6An7h4aAXS2CE0buTOVxM4NnhWzsNogZWYy6oUJDPq0gr9ZqusxzyfvXlOAp6OFAj
8hu+TuchHthS+KSDokomy/hvGuDmupPcuFmrX41HrAEtQTaBhpyBdfI8eG3hqGmR3Nh2zrb3KNJX
DI2qEfbeCQTXl2e3pVMjrS5B1Pp/x11QqtZnsKCXW+hr5i8xPW4LxGxo1WfMskVJ389RgcyLHCRI
3L4KAsw2PpSAkMzxa+GKr4NXh5Cso2A+nQIR/ea6WiiTmnMEqGsuxrSqfQf2vMIxScgmjIWy3pjm
6Cdn+Fyduws2K7UlZ2vWhvYQIpW8Gko44788SYpT9vlgTDsbheZxB1J93UBlcIOpoPt14OPMSbk0
mPfe3Qs51qEGnbtWH8YGHzSOyPGkDMiCP2wNqaYxwA7gJZPHOn6eiMpekORjG0ywxjfhD8Vxg9Sf
12HCcKmcFxGPlKHZa6uXXtjy55UZQ+jlsmRUa1Y/fnLXN7G/vETSVUKiA8U3KR2Mq4AZ68KpSWss
2d/Bb5VCExItVXbSakGIicUt1uP+mEGVZ/SF7TohgUk5J5yV6UXuNMM5ItiZfVWzw9plcMnBhNQr
AYZfa1TL76Vl77IHPnZsjp1cFMdKyY9Aq6P5jgV+IdaLXT7y3SkUV6pXssvBQI7yGgJDm2U/2GtB
GY2DcEcala530RrDDHN1EwpN/Pfa9b9yjsT55XUZUowbWBSc4dAFnTJyFGj1pM8ys9Es8jRhi+HX
lMC1ckX4ahbtckur+rxaq1nlEj8Xul/+Zha+2mQSpZii6KlvmiaOcJ8YVG1q4H8AJ0OVm5e1QAPU
ZQAN/9hPGRcgZ9dIiCB2Mmkbb8i6KHFhXOyYeV95DKSiaqn7M7kevSjnZpRldBXGIrBhgWE5sFpe
4wAP2EBZUeS41b3WWa30TRN58TrmUGcTGhHMSOw2kVmGiRt2taJCap/N4dWjZhTj3dABt2YQKLRh
FNXx5YZh6LXkaXijdwQfqywc0iCtqF+3gqeTTSRDiMGZxL0JO/DWZtWgxO+Udrgakdzw44+EzIXo
9qRD1nyPPS2M2ICtpFtnUD7yeQknNYeGCPy1QmuUQx/kOfGTK09/+H2u6uDTl4SeMm5TBz3Pb9kP
PigOX1uY/SWaAKjkyGJRr/Low6mrj1A6HYNv3FOexImFoZFwbcdr3oyPGkZUhahQIAVezR3rwUFQ
w7VKy6Ax7enz6yji5dAyJ+Tv1PY9fv+Y4cteMZQzuJggx//fHMlK7xH1kySKodsWDWsWSJmCiODK
qkhEZBWgc+8yXU6O2husv5Gs+7Cqx6hHzAHWWTPriLm/b+sntW71AlVsP50Azyin7e7TUnjM2fgr
E1m33vB8LkAkb790j7oRpAp7zltvWn8WNDIXR1qX3Vwa4vYGMmsVjXMzR81th/sqAg58D1+tyjXq
xeX3Eun/sxYVpLPW7+Xem2gQwnvKgftSxq6LM43DRuezcR2f0AueUn99+3/X5etHT21ZDpHKazKn
lPdI2eX7+JDRf+Qdqd7z0hJpFEp0Z02qJkcyUxTxOSsIXvudkNZ4+/TUeuabuxe0Nhk8UsjXcUbZ
Ce8dq0dUwbVdBMgAutpCaZCnJoHL5Xv103SYE7e00SWdv0EzxNnRwVTmUcnFs1ybZqzDDhdOdem6
3MmGUyh9+AmZUpDyLxxRTnK+jJXPffEUZ4lbKDU/SqIS4ggWVsnSCwCB8EotiHW4c9QelWvE/nNS
+bWjNycRDPDgbH49qBgjutXOJCDZxqt8yshnNw5ndG2iU/XrrvIpJufDPoYFRJvKuICj/y/4dnmn
TQQ53FtBmRydsNjcNF04DQpPtKCA39m2XpM3+Tg7sI1ftIjZPKeGrcsSM85EPf93auHyj7zpBKFb
+K/h1aZYrVLloihKi6gKYlNWho2s+FiOQfyvakAu/D+/QAbpCi5jkKJwl7vqiZos41TXb1J4SdFc
9aYC2mwpJ4VUJns4J4lkM2AvbMf8G61eFeaeKgyJXoetn4ypYpmQNGJIfYCGooPdpRrj5nLU1ztH
YNLgXnUtbvz7bUS5KMpsxWzzPBBD/LxYfXrQ3dhygQeZZ0Bwfnn02ZPyYOe4e/34VC8HGBp1tNGl
I9wRca12oyzDc9dieB0kaJbq/KLUqwACrxQ5BC4RwvS5hFyj8GiMDCrbs8MgIWXgWiWF+TkCbnuz
vocellh8/hZq0bjHb0PNv1yaCAIRDA//hE8uahOuHqJ5JGhLxdQux1HPjk6HZBXzaSKCONTeZk+t
pczg5+LAtVMjO5/A+DYffKZPacW4f7Rta+xTSQPGsVeOUPTM+1BXd/OMa8aMGjd3iYtZnkewxtXZ
v63huAje4rlchLIijO68M9MmVGkmGsuNIHiLNr90m9RNIAGNcWW5IaIaVydybjltQHQYZjYT7hOu
YUAZXuQri21mCksEuCLaoLb3qVrU33ECP8IYyzE5RuUAs2ZoFmL8KWmraK6pTRm/5Fm88G+JswDX
gXukCc1a1adbCJNJQ03Of5QSO1Iah92WR45UVQgKWlyu0kQPp/CDidk0OtFquDhQP3/jQRYbuNXG
kP4hwFVsPIenskLkZxtaa2ky5RvEyI5Z0levL0tfRY7TvtHR91MtHYbLOZCwQ3LnUa7NxaYQQ8QP
y/GrIPGqgnJSgvUWWOztWh95XSVPOmFRiXEV9nOwRivizHmaghUhJ2hYlgqQmiIbF0NO6rbHd/PA
1IYPivavHWoQFzZQLBHUT0lx5guXwfcmWhjdVvaTecRjATBQHYZ1JwFSfInRHVkyVOL7QgR56hcU
mjiyftBrB/Xpnm2wzBUSfK/haBTHvR0ZuGxrLkb2gaV8YEATdmBmDI5WlXcKa4pICxVPz1TsZkf+
VTY0VkTma58U4k5cxft1vpffVB6gBNsdRDPlPTIrCtDvgn4CyAzeR1K/HPLhOKqZWxGInoIssTYa
9S+4Gk2WhpYzqQF20ym5ceqjGwIClboab68HYPK52i/H9p4YOjVOp0xTsA9riyQIlCbwncnVqXwp
IQPGDy6wkSkkfGUKpBaE1fBg/AvKa6lgQrn3FVOqXkIS1+Pvtd5/kVe7tJ0s5AD1jmtNCX9KK1Bu
5pNNoRCokiOqlo6JoIrsUTNO31P5+w4JKDkUN4yVNHmblmHgfFKZM+mKKTjKYiUwa6k6O2I1AJvu
YhRSIH9ibvgE6eakYING0vbjZlQL4wtWLQEpKWLCnHOgxOPIjN309Z7Pm1Q7Aj3fPR3yXo3zAxls
Jq82ntFHjbkpJB34o+W0xDh7P6g78ZQGIXOhjue4WTMRnJopBgveQ8wARmxTnYqkkx5uXKugGFkh
J49KOVGFDvOOlcdcE9dbzBapsBLeVEgycK6GSeqDO3YZMFpYKCJgZ7r/j3SYsYYxohRadfCGTA5l
1Sq/uQUsiTXpvi1wmDN+aGfoFBxp2ltni6suBhH7bGFvwmY+F6M3DufvGwMDxvzmJzLD2R/lpPt7
FzU3CX4kDgCvDxt3SN1ZoKfQ/mVFpSc1owfNkP7RFMcGQekFHL9I6rBLWW8I5csrxPLqEfcFGKyI
Cx9dLoclY+Oym9eGFtodsbJdAmsGoXIFin20LC5ebiM/esw/nPgMuhn4xjUp9OJGHSfs1KVdtxTh
fN7U1P7ZOO6U18wVyou+OJFXInhRcQHDOKAE7N6b7y7ALbQGWwIJUM1i8eOiC1fmxRpQ6M+7w0aV
iKU+Jv6nMs43PPCUE5wnkViMb2E+db8eyvWm37Pxxtxjup2uruX7DOPVxySxVs18jBfrmXGREji7
dLroDktghlT9zz4fAYaMgxOk1p1HwWFF/Dyse5/tA8ZE87N4Nn1aWIrtFcBL+LEAvGCTrXVD+KPa
tvqHflYIORuNeXM+IUJb2NsqJqmWfVC7UKNsYJQobbnChOwVQZZSBrL3D1oT9cKGG2soAMJUFE4V
lncc1NQBFp8rBrMLEU4GyBQUr739r5/2FcA4J0Vb1HVgDG279W+GjLroZBLFgB7GPxperruyF6hK
IFGiskTYUR+jNDrVzg8I9e4EIMh1Bqa5RSC6LDhkGAx6pnEZ9WfUDD7zvrbZM2YXY75dBN0tbWSd
K7rqYXFQ3TZawQtG9ejByP40imA2ov52wbU6C6yj79DEpO0Mmu0IoiZelVPWOfAmbiTstsLuOHJG
Q7917vwTo2mCEOg0hirl9YmdJtkEDtfrKFWeh4iK/UhkSrqN5dTPHqHvEr9xRzatKvCyHw1YCePT
xsP1PFRJvzSPidfkCczYHMGo56+EuvhcuxvmyZ2UT0W3k2t2uijgLIhPC1kMlNiuquyy2+62lwZD
G98v4jke7XD1WNdz4Gi39R/uK4ffHrWs4vKJtbY5F0/y8F9BofRo8cEN3yEb0pj0p9ZbGDyGdouw
K0BiI9Xpld7/aVhY5hYADOey9HcJz/G8nSsflpm0qq6m2+FOyAxJka5iJlnuFBq7yrTzdFS/WrtD
7EmqR3/uRJdT5teV2nYR6eqXpPF6V5eK1ZDtxpS860Vwd6B1NQ2ai/PQ/WrCbRndfa8xJK79K6NC
FH1GntfX5FI2bqlZvmoj99ZU07G+JKtC/JR3DQH/V1StjOQNTI+T0M4NMJpp5yJCXVPA+1P+mdqm
XkihTL3kLT+Qq4D2BK8pIZdDx0laixLDDwuk7cstvD+3Eg7CrJ3ecFxU900hz49sbzEFMccUGfSK
ZMnP98Otojp2KR7y82v9awBawVw4Sl6fbZ95GbFmMaOISK77qyVvYIcbL4aqJN0DuzJjdRDju7Rf
KuCH1diExN8XF1F7wBecF3mEDkBwO7ICFwuu1A+L/oQeJvNOmOetmOgu0CWSmKSnJtL6iT1HcLy3
ScbnKq6rJygCApAtJXF+x+Wa8Qw/2IhbMCzcgJIP2DQml3VFPHV1CL/p7/fJpwtsyBuxWX2ddSKs
jDSpV7yStKpje68m4OFaEU7TyTK1U5VzJsE8dLVw4p0O0oMLgqza/K63h48z3beoUyEqhZEHg365
xodBHYMvM6vrv25yiIx5sAqlweq5j6gPyqJiltENFg5orVcBpUedFPm0sGM6ORNtRqpR3FEwItBf
JsOmY7NLAXQ4WJNCpgIegYs5uNxGelJeWMe9svLXLrwRNipBaG9ZtG/K7cXnyDQnUQ2g44DKR2DD
mNNw7zaDZw6xjf7aYNmZ3ryoMNM0THdT9HRkHdY0Pb35TQBEV82UQzDDOrV3E7DqRXaRRImYsTQm
3CCrzCC3z8sCJxze/8qxeXYCI4FdFh21gVszXvDjs0/7evZeL76400QTSP2C21G3fl4A0llmQ/bS
GmoklF0q01tJRMTakQlpQsM8Fv6lRb7OWWVsYJap4Xe2Sd8pxZd54e5z1u55oEiP2hVc/Wqixy34
iXHy9korLcp8W276N59rAewkJBZP2nYjGK74MTaBOTrvi1yWHWHfpfjwYPoGq4oNkoKPKO89XH+u
tIs0ZyqeX4YFz4mVtAXXiiJp9+biz6T+BnVgRMZF2VFjBu+EKfD2RErqVtIRks6RYFF72joOMswH
NKBlY3fVmzFG7fAC9D2Hr3NBucwGlGSQ+8TUoZPWQAoY4qoi7rTqAqB8Sq8Fs5swrykCq4hdC/aO
4WkzZKoS5MjfEAaGtnrqIqO0G/z4zDuGd/tCpKyTNIg9s5OkhtUKdrbhIHiU5cl9rhdHPkz2ElgS
a8lwysFv5xm640gDSMWiinMeE3204WCz1+x2VlQMDOSSYLL1CFJWSb59U4Dil7it5dVaKP6yT1DU
EVf/MznWA9DUjGNTbryi3mAUB5weDDFa4aBNcVAmQTGctaqV8Yftpb8DeLNGa7dhcCjth06sTzW/
Gun1ZT+7lcyOJly2lo5PS6jIJDZe21k/Hd1ojKnyqNmD7KdjOR4LW1qZ2KC0PViTBAzB3zdNFixR
1NNRcY9hzTDJUlID1cJ3SmPpojIJglJCOoNYgZ51Ae9oH0JK336NiNuf1NjTt4x+G6d5yctPbCU5
tyx+ZTEmMKb7gUJ2ChXcYi/hmFk+Shene96191IdKiFc7q9Hhht+JecNMKSNNNycXQxUASDxuQKz
KDGPzIBV09kbl5lGfLMg4VlMrKUfJYrGz3bmU9c1vYJ0t2azhBxi4SzD9S2RKFrKAOYOIWDAEyrv
GEUWsMpTg4a1q8CpAj5fhdXiDMaC+CmzqIhb/m0bqn4hIc4zaLgclPAMs/lo+3KuA+r8DY1h8u5l
4qPgIv0txMewA/+Y/dOhXkkfOO7mEycqi3e7A+Zl4WuqEzOFne8zhE+Tk/Ni0hL8YE0JGx8KOoEs
BeQbvgWpLLCttRISjhT9ZgUujw7D5N4sB0XE2WovD0Yi2WszRzdDuwq0nvaew+6QEcVY20h7kwWy
HFRd+ynGbZWDLS6/15CoSQ1o1JpGhOaMm8YRay+mCHeip0wvrmQuC1nn2s6Ytyc2Odx/bOV5y3lL
nTPkeQcF5pmsnhU96xygEjBlh9RthiY1COmXXWqerUIRmx+jsDzpL1d191uJyPQz102BpRw5TpWa
wlZUDZNUjUCSkEkWTAdBaK/y9slh24DyTx9KKc+4c/Iiq+d16YulOebq9C7Wc3E44sRU/fL66DQ4
l8z2XfIGz3HE4/UEtOyyzE6QEkQb4Lka2Ggnxf7RxQAoBSlOUCcqYVjB/jJUgYeB5BzTou+UNHTA
H1YmFy3X88+edMmurR/fkfP3waTXrnrjoBoS5EZZApoWW9yxtW0pXgBoikAZ2YqUODkdifdQY4l0
FjKQYPHzJF/aGRoDREHfIAO8DjZBhhlzlINMuy5srtLrkWGBDqUFY9Sp/MWGt2KkzYo39WxyvKbC
iDuv49MNWCsXnvi4KcmR6i0c98jcJAX/3AqretaKcgEisJQPkNHzIW6Ju96DhOvIJXpLpbmp05dU
7tgujfrH+vXINV5RdBsf1CD3c73MY0+Gx2FuwjprbZgLwxGRNVnrvP5NoW77U4sn2CxvOXSu+NF4
z+AT5vW9crxdSjU78LN5HL/u3n6MoYZUx/Lfc/DJs+erlG1gJGCDZYfY+h3NmKz8ih9bVGWyBUpB
E3Mnv7BFAOvF1DFlI27rBPAwBoBifzSpYWg8xrPODxwMMXxlRdR0JQ/cSoy/1BX5WRSOfwfi6TIo
EZV47bLdr9uQiPHrp/W6xJrE2sGYa8T1Ju1GhvG17aWmnz+EU2KNGvvkqFv04Tm3BTdXd2G5TWKr
3Vlm6iWguQoCS40oLRF5bTZh6UMS7hEzTzv7uAQbDh63DqlNyMoq/DKbfC+axsdzS8lWSdRiwem+
flZbDd+B8EOm4qxtmj07sr7SZLVh3b4E4K+B6tYxtjKBKQnqECk6CeeWusKw76vQOZTvjbdUg9VM
J4uYMRstchdiiHEyfV4Zr/4DbitkWpjreb1QwYOEQphBQb76F0BFksxFZYQnuUoOnnlGdVPZOhyz
5pUHc71S4F/FqJW39/g6uz18Oe6A7uavJenvrhp2T4CQuAKNA9t4GNcgJDCZfyU0hz3Rnwim1i3+
haNziDcZsK8F2ll6ijHI/pooHmdj9ve7gHrKr2F1D3xm318u6+Pl3609ncF09CLipyVZ1/LjJMwQ
nNGEVd/AAyRTh4dqHrKNw2e0xnEuAKFF/rD1SMQ/wxtQfubJHEV5Zq65S4F3Z8H8BGiTm1nJ5djg
a5cAUdGyJtvOkaeKpa4uY88QsO1A6l1LEhE5JK3sHVtBp7zF1pB+y5tWfLYjiYrThazmLXInF0gC
HipoTLDNSPrI+vvLYBqmWIXKHdSBU3OR+LqtSwVaAuk8AUBBph7hpPcwNgv5FT7UyyrKBMVtLyjq
OOBiI5/zlblanEpss7SkbES26NNp0sm/ycqcQt81okEX9DRbuonpHxAk21BcykN/p//Nf+YjXyUo
6oaPpuV5RSqXHsXw4VhKZvZHBFWUjc5bBbMEBKh587z+adkaFD7ls2yKLqJohTYzfSTiRM0XNAQT
bVWWMly5dsDWVKGTDlO0E4+xanAFgxa9UUH+hmdYf3PU8dtAS54h0rQAlxBqr72PVppKtwttok7H
Dx/dXVfbJzGXGJp1Z+s4Q31HAV71b1SdbrGM+nqEjKkbTcVGe454RrKBoeuBcSfZfhna6x/60aX2
zsapfBuoncbPCzJIiSVBvbqUJ4GNKH7VgLMEKxpcEf2GFaZWLTPOAN308wbyyrKBD5vKnI/NDSj8
vGP0nqR5u7xG/1hHUD+QUya7SPZI434mWTsYEgPFTiO7e5Z9EJVtNnn2pOs4CKAtES05hPCtwui9
8wf0c2Nqc9IuuPF8rCUU0yf8/FXF1vNfXeTTYf/b9He8JNgATPaN2qC52VHaEu3MQGZh5DshkRqm
a39bJc0ob7JMTFLCrV9R3gC0WkmUMI62hC01trN1ZMZeVbOn1StK7cADYnZPikFP81sVnc3+RDde
j+SYuj8vFHwtmhFLL0haWc24UMDGB2dkbYvYs5WmPd4eUnAzUAm4FLaGF5TDpXHN65yRAXOmVUNU
LN46VxM36ZneVrK0ilxI6eVF+RiWreyap8WLW3uLSVq+Dv1p3O0wedhW2hmPRpkELQmngH+HyxlI
aTauBuCTQ/a35mAS94565PB0tK2wXnTPG+JlDTb3C1JJ7dOpCasd3iarfVl1wQBzFtMNo7xSPzYu
nsQXza2OtYiOxhrUY/s0hBCq3HWCeHdvgFBYtbdB33evWxT7OuLiahGrY0DrC94BhIuAf65/rfDk
1/Bo6lTgSWkQZ+SzrnxXhxz/beTs3apiVRC2OrFFWv2E/YjMMtHnVpRUrhIdTzBnxpWUhKvhPlU5
bv8ae4pD2/Ak9NzQ9p2Z5Vjetcbl0iH3X8Jn6JvwcO1O1C2gxctpn25X/ByO0V5x/EbhIvLAWk6E
m6NzkkFkuY8se4a8IX1GuEjcQ44GgZfKRU4zYUFwozX5xLvfKD0Wx5r3gwvix8UXq75zS4FGExty
TyhfnvPP2WJ3uzbvat4iT+SWmQ6CDNH7ZKSGM+VUphudfzuv6cmIpGPcdyV1+d4KsYckm+j8hd8t
mCeag5J289Yo77gSFlDMPRwoMOfXEsUZ/0MqsFhHOjNOL8U9YHwSLLA0kTrm2VXm4u+bDpus82yR
9jzYxkye4R4R/kkuCvcRJtlvryMIvEc67itXXmhZ5wzjDCvefO40s+DDbuO1S+foFhhaY04Sk09c
Mh3wITnDM9SowXD18t8s70NMJkJD1R8SsdiI5KAkW+4eX1QQ6U0ZrPjZOr93JjcC3/35oYteYjI4
D31+w7s2onMFjF+E8nTLh0csbnsfH1xmWzVsEsVgnDe6iOaYUyDX/T6cKgWJQghpfMLnz2BTKrvu
E2IQZOOLRjks1Phop6seV2QZs4S/AL9Bt/lSa6s0lYzVNzggYGFHXB35iVfCycmNq5NTdjfzCrkd
Rho97Djd34wYf0D22Y1xSRwz/nkEsPZu3+BAVTH9D50h+gYlsdO1Zj/5tV93teZR5Zw42yfugKJr
IKkO1Z1D3BgKGaVLkFh8FUR3gM8cAkh/u9vlgHLS1YeocuaTsJgv8d2BiyuZCBS3OymA0MWv99RI
UjX+8RBRONmwSFmRabpiPhH0VDiA9K6oZ2ABygWMEnh6t6YNGQGLIqYOM/UDMFiRCaZNc2vNPSa8
A4gY7iJboofHcVgjCmYekogZMv+i5H5PPFCWFO5uckfic6HEMF3zhvVD5Wk0cE97diWTSM9bpPeQ
bJYkK6r4jGIk14KmpWP+n7JwdP/VIqwJjSgb65xh2En1ebcsd1fg5giGJgkGEZAU4ilNM2vzZxR+
IKJXwROmWE8hCVYzM2/4lT1UNoosv54d5HStdlGD531SqvJbYoPcBXEksD6KcFRpTMqV3YFWHsUJ
s1E4DqUUiGUSZTShhMw7VAoYsLBGOsdb6SOqrct2Xs53z6I0yEF+ZdcP6H9Z9I9WL3i20cRvBboU
P7XS/RJ4RzKQKjycLefjb5JNjUtZ3FWosIg9kxDBMmgBh5YFoVzcaY3qU+/rVS6R9+f1X4kevQWG
Y3vS15MyYEulGB05Z23btlKbCFCYPEKFHOgTsK6VPdT5E/lZWLU+9uwb2eeZ60J4p0f6ybR67zWo
57XfMdbl9ZWYM01aAJ57XGpz5M8XdE1knm0Y0VlJbiQlihiUhsbFHmbEsNM/KwesqRGV1ph+Li58
3ge5uxYlzBh2U66AZcVXtDFitOCJ3/vMZIbA+XgMw8y38gX7/eECtS7rU36uXdLxaT/lk3CJyuX4
J3PqiZRLbNjBXLdAMTm+OHcE8XHRLV4bV+w9n6m7EuFPCta2NkPRr3FBttGmwweJBLZHExI2ViHI
R8e/GdJ45ndxmQCDdcQsmZCcamyikpEaT+kq+Gs4Bm0Gef20ajK5mxBsjv94KTodNFhuMl394l30
wufJAV//ntkfuzl2HVf+j+qoDbsF3qCbhoWxyq8vwr0VsAsuMKW3LZ09qdAzzSI1VOfxJnwkX1b8
1SnyOxvsrS1yVSH60d92OiDjQlwzxbVxtUbUh6UXMCXQ9+pBdlWTdt8jUwZ0EFypo9OR0iLYOlDl
RpPhKBNJMX3ywyQ2fzNCRPynOVjX/klk9rmGpdSjrbAa4TmZ9NMC8h5n0L1pq+Nz2s88H56D/6q4
KdE7hMEgV9xHbdX2E7cvMEr22zBorqQTA3u1n3SmAOFCEVUfCMbG0yk/WOXgtE9FAnYr2Q1zCRyD
SREvmsP1vd9ljrXv2D51TV55lcuzcr46D2RRHGObs3p8eS/Tj96r++7us2d6LstCiVhuejUNjZ8B
UpwGePSYaWYkwVCPoJ8kPklFTws/hSTubWifNRLf5Ll4Itb6RN8mUNkI3I5Q1EB6ooDMrIqucFOB
QSvd2CSKw8zcuOWcETK0OB4oZHvje+UIXbWxhLr4XnqVUhI/zvYYQAyqnaoZkgsNDv8rXGnl+87D
Ie0mWfrIQrnutgY/NVz5OBvOEZZ7eva7CHER1hg0wUWVaW7iiVY3oAMBY255qkXNLUBaiF0e2a4K
TP9QdfkuGHPlxsd52Rg4osO5JXVYetcaG0NBLt9Z8iSHbnteWMAnmPrnbG2YpX66DWVIxNA81D1q
tsQlV+knLJS6LJmmSod2THOMcCgNfTjsXWmoDBjjPEca62Ro3OjaASIWB6Ba5nBAlf+XNqkIunuq
NAJwy7DQLCqqmzmE7Ip3LSZqWbs5nh2+Gnm55eA3Ys9f2ZyOygmQ/dnmXfw54LFdnLXFmWAFAee0
TNgR8PObTELe4w5KdKDUChhN6vvZXnDf2GpcD6XRy7XCXOD+rwXsf7doaX8ytcIoP4q4gFIT5VpW
sJcDP4YbvxxdwMz1MYP6lWkCDRh8vbRB3MvgWAHY0YLoT+R/4QN90cliVpcdXJxTM9rGHm4XWQ3R
DAB3SGK5GtfaPk2JDGUlvhaZ4QnrI1crb18nZUel28NUXVHDARjSQ7ESDTryYTA7Iiv9GVPc2gS9
lnG5IFbs4G2x81/PuI9RwV7r7PWXg/kuDu8WP1GMoLd7yl4hl+chYqvn3TT0BUCxNByj2TZXOSxK
wXNU7WqtXq2f0f1D0oGPr6e5hiTKAwaa0+o4NdmDdG3vo43ke23nOYdJTH5TBFZXbQIL+ChWQTS7
iX9L6V2LTGpkb62irdpVdF93GTNG6tZpyAolWfRDiOhnfmQiMNB7N3y9KodkC5Kyvblj+qSlcGXf
L0E6MmmcM34DyhIi0mtxEZ/3ZaVPMgJ8nn/aO8hz4AJKQJtFhBynnGbrPMc5sWS5LCwjZ57DnwYC
gLV3fkFT/QNVRzvM2yaiWUxc3Kmv9EjMpYFj7eDKe/RbvkX4FsDHKgxHsdZ47GCOFA34QA40ZJ7u
WElGJj4mH3vxhz/uudspLF97WnvnyehZI3NLZdeh+tGDkTG2jvap7EsQxmoZKcgmxN5B1ZJqM5f1
vTwM9qc6Ur74LkzFrcx/+xtbcAeXkptD8eaYACJq9+Oqotw4a7VQID6M64hf8Y9F5ko6RqvWk2td
F+klpR/MrdLJcbHrin78sa4YYSIJQ/MfWGeqbf+UtwhYCnRUvKBfs3MXi6qfWd95o3kqm1C+hf36
Mlr7U6WXqg6Te+1/xd138EfxnKGFq+EoWPuuF8sdDxkhXaxIh8E50upgrV0B/AU8E8N9dLewpBV9
0NXm/0y49vDK/OH1UheFs8X6UzXYfrSRjCy6OrUpNfTYX2Q3zMugbkuKRSdgVoi1RCTPufzimogs
F3kRfEu7uhe0ADvLOAXq/Zv97XO8lK7X0kCczmTJvEqCiKXotzaA/ZfW1OWpixeoFNaOySph4Lmb
RoS9kOsJitB0rPYoW2j6jV5A8lMpS7L3OVB3OZOTIj0BP890NUSC7fzQmocBH9XhAvm03UEaj7E3
hA/dWGDlElLyoPpeh5+dCjPRkq8GeaEokX+H4VEbDjUtl0PVRVTOwAERw6isPArIflZP+KqyXOcH
2x/GKLaEsUgVgdSwA34BoE5YMTO2A0j78B0ybGKBYmezCzyNzWxA3IIJs4bhUp6AxDku9tINfKOW
rPrnIR/baYeBtnLAqkKT0IAYMwncZZgjG6yC+HoODu7w7NlA24AomTUQ/qc724QxnGD2EQ7thoox
Cxl2hc0zmMNRJHwgZw2iZUzRl/zmX0n0TBvS0LVQpa+pBlnBtli4IZ4wln4fsK9JPTCLad+P8+t9
0AaFa584a3pF9tCQAiefDSJDbiNzPLMZzvxl2Aq717PNz10R3MN1CxAVd81RkJk0crNy39c5wOo8
ewENj/R7sB36fZHKM4/BtkhVf1uQNrx8tWLTfNSJ/e8VoOReEbXYQS4fHGEaU9tSd5cDqFjjSSEx
+2yC9XsiPbniIGCg8jTVCll+2c39wlJQF6NBYNnYV0De7lytXAXTj1mYCTgD6Uavad3zRLfWHXp6
FV8AkoJG+zcuLjuxcm505fEDSDSPMhDDQWGwlJwLpNr7p7SBmaHn3vMPlYu1NfRs+/V2EqdJTVjR
fj36jr08wfHDoFN4icHY0IQWapwoiYgzxeJJpeZW15934ioltcvuy3Yc6c5QtE0OT2nqRmM44mB8
OwrV03ii2kunuXzyTcZjlZjCXZQyYvkQ57jv/klnqa3dEUgixPvjZYkSOgJftSgMPXc2HCr6ErXQ
Vb/UN0cOXAwkJCPc9AY6WdKRko0aX1G1ddL9WmUok+a8bP+QlPypNAu4KeSTT5ntThL20w9Ct2RD
OhN2wcvFQvsSeuYWIn1lT1F29ZOGzOtVcq5Y7daxJuu69gbVW8WTRvTf3hUa12oLvXW+PmuizVpr
tKFeQHgfoFf4GWSlFNsAb1/N2dDxn7EzQwIvKEfWsSNiR0TM411ZDqKs4+mKUvcSNAjyiBaoSDyG
AiHnvv4iN1P95vhix5s6dyii4QBrRSco7/aqdmuufZaz/Chi78uW0Z8muhdnlK7oMIbSjdarmLXg
X4MclPoC5/OyXOfd85FqsmxqOMN7F3hbWPtOtsT1md65+ZV0f3/G152Ti0L/xFsu/0oFieLMsSQL
ADC1iUlnBWloYVqoI7+dIOvozd8e/zDo/DFjzvzYcXv/tJUtj4NZJAjSDFRwkWjzLA8q29bi3RTZ
SzQrK5jNuS0OigyMzXXUm2m3cFKbxoeJz9fNvBt55U4IPUVPq56GTCzalszN/ViPGHj3J3ZxjrlR
6RMdF6m98qfnTDUiotEWtcvGPAs/bqrV+HCVCBiQIX7j3iM3h+zm9gZSGmhAyoJB03lYiJ7Ik37L
UU+4+YQu3FrF0fkIxVBy0uQLQzh+AJer6yuRwmdg12wqzgjpLy6CXKq3PSVlZYpcGVOZkkPHS5HZ
72Jj5oFFoHj4EsEO1GULEbnVqQP+W43VGJ3+BLWqIFJWxyi6tIJhvU7FyD5VMs1addTwUUr4PKcD
6nW9SMdpnpkC03KtBGTjiU1NhWhr36eOk9aiTCq6VEzYsFsVNHGkldDbsf5ABUhSj1UEr0PM1zlO
fK7DPMKM8/BwkV20PTctqjfuNpr8Z9M/PKnuHzUc65QsHaX3noWUuqobufPOW63yU1WE9U1p3HTS
sWd8PfNUGgWOgawjJOVfypCXBjMd2TIZvt1WaUy5Zxd3sbN0nmG1ESQ7waJNM79TBbWf9vah7f2T
q35WRPH3PyADbnKeOhio6TN/D1dDoqtCLZ4e6F4Fj7/O1su75m5W60dwLM3aSMVhstPjJ5Xuc3PP
hw/xWVzsO4yxkv44HDW6LKpAFTapPwHZmp2CtHEnVEhWMNeCmvav8YZrvmjBvVpb1lk52Pcl0JQK
1tVgAE/hItRY2ncnbDfXNzRDR6NYWqFGc4yHCF7N5u932o/8NzmHdyoV84rRaUzXAiSmTAAypKqd
fpE63B26MmnZpxoww5MC+i4FSpaJ9UOq+Tz5QAL9tyP3IyjFd4ZfsCr7xbc8zXCqHmWf9Wzq6YbA
xdTyJHbVGNoU0AZfv8bIqt6DAB0oTBPDyy5vAKf2XuGl0UbTn+k9+P59GpwRJOQQmUOyEIIeeYE+
gZepY6y8Pxm6FMbPhtxevCkX2yTTDj6R88l4Yp8e3I1QqrKDrIwkbfcPtrGyHj76tK5dd833H4ZY
W2ciSQKmKk9YkTWS1u92jpK7TtG1vyiXaQzq3/DFixDMdKH08fudBX/YGZnE4JHQcel8tU7RgyI9
prK6i5hVHx0PhLQuLasEY5mBeFzh/TpV6NV5mzaOUmka6FXWEezTZvKhCALUMjY4orFTbjdBMVhA
dv5Dl7salq/pWSnScGOIXbyGMU1nKKjdhSubeLMhYFhkZHtnx6ozR6cqvLCTSSdMCu4iox0XboXl
xPNmG7TtOYBoM1iav3Tbbkpu95qRAU3C0nIEdxD21RVfE/KwK7hV4muSJamvHJ263LpdYle5Iizk
0ug5lTroO3gEeClcx5cRp0lpFVXD16YChRPP/sV87bLOVPBKvzTLp4sJRYwQx4LQUULEGjXUeE4q
O44mnQqkSCgwEsMM1VRrQudNnRMhrGtSPT2zrKOagb+ulnK96gYtn8Gu3HdWXIiUTj29oX/zpInL
Q3Q6iB0vKvdqVOE3dGL1QQ2IcNrI0J7xG533qth2J/nyIyQ3AlO/pBDohecMz9AsfyG8jaij7hDl
97FEm6a555skz6B+rOma5JYHxZOCwv97JdFp0XZtgLEe2exGQTlRocJ06qbNRpx1hW3d6OQkDCQu
V/f8j/4bBYOJGArpTget8ktCWGj5DrG7Nd5Q7KD7j/58nkU9ti+nVGjPxUJbn5i9cHsofD8OkxoY
XaG4L/kQ/SZZvqlHgOKZkVT5bIcQIR3+d83RsZOvJcV55p+f5eqgp5YQCijC05H1OcSXlY3Mx4fD
BNMFVCkYl9TJeg+xrnImezTRVq4myCFGvW+jbhx//CJfOV2Yqbn45cg7anMUFGnvAdvmD4S3qmct
rYW0q5mVfoHQTdBmq0HrHMQ+zZVMSCirRqG5OzfPGwHDYbM0kSfQPPoDH64CF/AmQHpPyfB12HFT
Fn4p0omaZJlCLAvoR8oD2fW61EeJ1mqjlx+B9aqkjuaLeW0TIounB6YL4vnFJPiOend4pSnRds80
bT7H2G5nntor5AcYsTfNBFPtVsnGLnn0p8YCgsvkbvrb+6pERBf7qVE8bOWyyRrHvPkqxYzrAfMU
i+3VWGuNORPWK1ounUWWZrflaXYNzQALvIEiCeIAxT/cnzlyCuJ6tj3sXAkhg10BjB/hIuihYNlv
UBh7UE0zFT4AniMyD2BtCDRSS/JxsP5wge97Hya5mjGq8UQ4//81dCbUBl9+tIyxt7qrEP8SEe0e
4dL8wDhmEnNrqOGrSMmWF5O5+s1pOtRIEuXD92wZwYSiYaGjXArySsxrMiNjSNXN9pM5vtFKc+Gz
CICtU9Y0jfdI7/uMRok67wQBN0i0m0BdNd5U9pChPC8YnCgCGltyMj2nkI7unPJNY1nphDeYBPTB
QJ5oljtZ3Se6A1fhUrSU2DCJm4vUckz4VbJom+eNd1Lo/NdrlVjI2q/KExAdN8EO3WMFfsRNEyOY
VYc5YSpZ2xXL3Xcvo3pTd/zj9VN9mRufG2Bl1TiUQqRfSnM1JeMboQ1c9yuXJvk9vwjPvr+2gxNG
zqVxG+y4hnwOXPlANxFRNuHB/BY9oz8LDOvTUA14MDZysOnPgUHyaf1rKh7DHUWKWg8tJoc/9um2
4q18IN7+NHzK1TxvEb8AQXvTcq28e8pAi6ky4vMKYX/yxZHyeBxx8ueJ0zr0uNvTaDQr7yma4JoF
MVV127BT/3zNDkG9QjOZTtxh1Fw0/LkM7smXUPKwWeekDnvMtWjwsM3jlTA/gX6btq+mQ6YK4Tew
7Vm0mSXswZOXvvNCUc0nU4LsXevL2DvdK3fdpvAk1LOlom3VM/q0mLWhSJdy80QLH09auJYuFOL/
DmRI3KDg+h845jc0WtTeD2TbTaynA4WKmWAfbiFfNlNQrqsOzjIdBLo3XWnEhuGff8aVFtbBuy4C
VtV7PMBCy4Sfg5EozCmNTQCpSxdvyubv9j3M3GpKwSSDOjNy+0SpbjdF/BxwVWOiwNYVR26nckdh
a4GIGDiR8vtB9spYQxpG31zIFvx6Drszjwv/+YKieRyeQjZk1gpRuF2Gp5H5RoFPRICMRMMOWHAl
fk8BKD/w2emtiAFkdaaPA7KaFS65aT3espVbi1lVrD0WJXg+XjpQBJSnBVfpBahINlWMYO7E+NB1
7+mAYH1lPdOu/mA89CAmosAQmDWQQGGQ5lJUpvHw0OzPQKWpZuZWu2XKlnemq5caYyfD88V9QRz2
AuAyJ4XlzuKQpz2WHbNUgurNqrKP5GXMNbKhd0j/NJfW1RDLLAWievXlYj0PpfPHMTMJ/SxVNOfM
l4gy5+40jCPn9/GDGZA+wTXyQefE6M0jSGkWS0duGzZVZad6s9Wav+UCauwkGQa5dg4ngD7Afmto
4hityP2YQcyXs1uZ/vMN5rA+cVQ71GIlBiHP/MkfTX5zQHz5/2aBLA/EARMR0CrITP7fl4uQBKvO
h4l2WUcsFLnnnA8oLcUU4K0cB76g8batwws8uR5TGhMxdDp6d565a/Vxq893UKPqsyKYiRJE8tQ0
6qusHY2ddAlXAaROi3OWhIQNr56jkWMjESUjoToiYdN5JagvO+7BB5TYiRXSZvnVV7isnN/6D8e6
uIm78AisjKOZ0J7RjagPx5PvwcpZ7hMlmD5dwjIVgYdc1X71fR7vY5gVSXhLRDL4IrpTNFas+oTq
45ot21X1u1NkYgHL0/7wT/CepGRTUkqX4Qcj3knJfrP/gzQWDLXYvRixmGbZk0ILTrqF1M4z7cZV
hH/hmaduGQwJAATYrsNPSZW/pu+RM6cAf41cLmDB7aqUf9UJzrio2vU+Ul2wudc4JgCUdengaEKB
HmhgG7x3YZltJxoWjL222VktBWrKxN8WHNz8I1Sfq5FvfZXKJYlYmu49Htuf9YpnM7MOxlngqJ22
DcX8imDA5dxin47Zn5Gk+phWIVQTjSXHwjdDVn3IxWLkBVsJznYyYSDp1sCXrBDuiC9cV0EKuk86
MRKpnhcoNwF0jeIv4EQx7IUQ+XaUg5awiXljfFIYD+a+pS4Kz5yza8vz592qSjHNYFXwHXxDPrkN
hgCsO8VLmcfO1w5jPiRVZL+/u9llkB2EQ4pRHzgFsoyt41AfLzAUzxdTee1n9hrudEwQqqV1XDSC
uqT8tL/5NXSbkd4FuuYM31IHWid5M9cC/TpwMXnUA3xuDMB+tYVgaDdmzq7MnD5a+dZY1m3slhgm
9VIBi+FCV+OcGbDXlIN4g3dQp3XORLqmSurnlBH3zCFUtjUUyC3uryBAVchZLW+3W2BblHzQM3H2
M9Vn2YvGH3TlxksBq07HXjhRZl1rowj05qAaRLwsEsGQMT8AVLRXDgESpt0YSNKyFRJgKqCJwFfK
xm54oLqNKujk5KshEFCWbXMXcbqLi+9g01ijQp8TRIPA2wMEaRR6WGnidI9BIj94K+sXqmX57lJa
FVa12YqpuYoUrV3Yy8hilTonemhGrVlSYJ5rrEOBy+QxgB9elpKFmHTu0bJUmgjPZyGPluVy8uv5
gdPTGfRgnUxG0FeSiEm5P29J5EIZSdwoNyoPCYmX5/xmyHVPUJHUPMEzAOUd3A2J8Bd0P8/8yMEl
H4OOWocFtSUGeuN+tUY5Y0KgSLTNOwfwfdhw7q4KMfpimWpNSTYfTV5m/z5MtMhYVY3G2N8Drfwd
bbcSOAqwQlKKu1NkUahgG1t+/0ra2JowQcsrLr4dh4hzDKfWevXvp1mvoNIbvOW8NOH4HE4BKvxc
Nhp3xVVdFoljC4Jz78P6BW6zN1eyfyr5BjmZgEladeOFHR/cybkMJjjJgCnuZHxCjjX0E//YsRki
Kwi57kDsp8BCveom0EvG5+Zg4VpbNYJX6W6x1bpZbFUhjrOCCXOkOfIV16M7Nu5e7+k7pot7tJ88
lCykVdFHEUyqjRviqE8lhDReUXMumqAmKA+lLqA5oEZ1Ld0BThgHS0kCqo+EL9LgZYw/gh8kAv77
wmjYf8GcKqitmTDr3S7vXysU2o0IWFb890pi8wl8M0ju+E0JW/3HTyuUrdjWokXS/c8pXxGMZ4zU
lwCqqNVkLmz4nmUnti4DkdVzykeIMZ569eKg6/S0+wTQKnRHO12a1qoANAAVlol9tfZi+VhZVrCg
MMOVaxdjar0dhz4TEISphtv1UrkKI9Bt1+JaUQPgKe76xjLdleNXVhQVb5xSRD8i5TGr4NDmdZ99
csd5m4eLu8iWPjijIcjmQQ/ILQmTJslTqvEAc7DalhTIXaPTMlNaUBKWsRjo/6c9M9vxXQbh78VX
0De8tE0fVYmbuPjiJwb5+TYkQUE6bApoPuQ1VwCDoY/XKUbK3IR240x/MXZdSb+Ch24hKokxNwLU
rO96jmfT3NZhwppepSWU2/d2FYju8kbyh7nM1Lj55tUvRZOY2X8yshdsWQAPuhzYtLO+ZST6AK9G
KWqJeE5m7q7hdsVAstOdE/Peav9PEVyoKmdIhtLKTOwuAyOk/jSJdm8RncQxMbW2LDeCZArafqLc
59kT8S6y7c33CcpiwNxwdktzNjSxPXFkGbIgjV1YMfL0vgO+z6UhbO4IQRMmC9aMrILGWIX2sKtE
k2q/N+nkcg+0d+1MVxg0+KdW5MTm7387SJ+/JLPUtxTxLUPwxEOgrKcvv4WapARBaf0pRH4JGwVt
Exn7FiGdlzSHBsu7r8QgmEI3dNQOCehwzNAb4VumFOCO2fiA9PDhkrqn8YAdYiq5M7jMez7pt0uO
uupi/IZ6vdKmaMw359ppSkioodxYBTj55gEZSvwXlMeXUxOkgoyJCAH+srsmP39a7+Hu2EDySlmV
drVS4nnwQICMf7ZBuoACV5C4Vt+TWGcqJZFh3cLf4m9wfkN9RKh7u6wji9d1DnKrqM0f31xccGfA
odTLbCABdVSPae9RMPF4aRXM7uQ63DMjDpQTjCw0tfKTtOCnoSUfN43qL/7cc3jA+/SfzX8elVaz
eHIKKBVpuMmy5KpAKYm5E4RWx+JXxfWtWPc2ofQ+d+6r35rPQHH1Gx0OeUMHyLhNdeZJDodYOKwr
VdtQJDWph0Sz6evTPym6r6w+u2KuEzC9VlmsXHMgca9p88UJwKuQLlfTBGizfwSHXEcncvr6coBK
BujZj6K+VgHUhsKi9Ake49EUJHLHp0eWK8iVMLifp3gmsg5jcCSOQ2bLJ+AQ2SZSNQr+DdZnJKZ8
zyup0ztFA9uNd4g2vcr4GrUEomH0VQtBECaF8JWD5f2d4HkI4kEpTlpdMb5uPmZiffF9ri8jGtuH
u0Z0t2rsbYQYTWwIo0IYgQ66jDHzVp6lPRH/n+yOJfC3mAc2qrd1BpqSVh1UwjepO3ew5nyiXDJC
ZbTN6db6foinn2o5TXtEzCAzg5mNHaeQKHSQm/5mEIzeH4W1WOvHQzE0CL2DdKOUIKgzt9s7UfGq
vyGe28vYC9HnG5//M8ZXcBgKOLg8UMfEuWqnS25IQO+epsmLMLnZdciwhZAQsglm2LfXMJ2iOVs1
XfZmRIXTk2ygMc74mEEYk/wYyi1oCi9A2hOj/KVzwEtcLxgWv3K20ReXwOqY/OGfss1uv8pFzWew
5Zw4uPLq3/ZaeAiaOT3gaqRC9M7p+CBfcPVxjtsAkOEUQ0jR9J/LjgoS2QvwtGPm2k2Tr8hDQq6o
YEBNjnipnvDD8idWyjk4kAMMZwb/e+JaZoB2SMKp0MFTfIs7p2V3CRenlHH+ohGcXtShtAIb8ce6
ED8gtP5aLjuTx8MpUPyfiNbm4u2LIKtu4P/5ruN+6LLAmxGU7o/rNXAr8qBeINuMz4fEny60YCOv
2heJt0uYb3JuAjOaeDhkDuW2iy8H4DN/t2Zb/J5TBDzZCDnkd4DUVX0l3JR7mAYuad0e60qXQg0h
IZac/U85Vn11bRsROVeWrjbXvslt85uHKRQaXfJcWA5mBCeGo2Gl/8NTlQWbkKtjkcfvbXqxW8CJ
emj84Sn5JCOC9xxnK/7XOivFrwQKSVTxGaV9VVOED/3LJvBjqH51OR09m/ZEwabtEKijjHWrRF49
vviJgElkyCzjCxwx2YTzje1GdroG1YMe/RJWZnXA0Gq9M7ptgePmieS9MbHdYGiqtnHcyz/vArMw
DOGDLO7KaCQI7XXMKEwfYSxTh/X8HC7rWAmZDEZtbsFxsJIKxSZprOyzzpKKLc7QrW940Wv+xWlw
NaSxRuHn1Oy5OMK0uTojLqhJLiqW8JT/+MU+uczwnIGcd+Oe1P3xvh8IV9j3rp5wQApYRWymegAa
xv04gDGTMKumGBO0/UAqKYtA2D/A4NWIwSwhCHejm9zP7Q+y8Rhu+kf8QAJL0zeCsFm2He/JZ2Go
pZKd4u07iu3Fi/9k+U/gV5Mdyc9G3tSXBN4A8/4oQ4+JiAxTvCu+d1hmopHQB2gl/yVer6Ud29UU
auisyhesMtoAkbDdnBvkNMz+gUnmGcl2TjbCCeBlXL7GNduan4ruTAzobk0ZoqqL70fe8fws5A5f
HFKB5PPN6r8r5mj9MfNHOBnQUE7y4jMADl4cUhO+A60mhsrMZOGmRoI06UFwyrGQpcA2RizDEkjV
KUtpUYttxE5kEyF/lRFcQS1tp9Jaj9RPdYBWAm2ZgU9CShXusOTtQZbbgaq6mGQydL8xpa6rG4ZF
/rGQKfImCw66yy6YYccX5Onu3ZEGnGmITRLFOvrDI0Qp+fZlhDK1UCZlfTq5c/GllCTaW7Q/O458
ZMH+qknRUmJ0x6hbSOQR2buhmhyLUxi4tUcyM7bOfmLWVenoT5fh6t5tq4zuK8oGgJPkqgwqRKoB
RmDtxshvILY3Ec84Rd50p4Fimxhq4zDsoXCnykbBSKDgLjjI9E1TA1wAWSd1qdW7AkvedH4bWuVz
SMGjGIlr7nzh9hyDcIR2zqLctdSjQx7TVZGVBqr+lSiTVwKEGGeFkF+BLSMsR3eGl+4BFqyR6Qoz
j9sKB+LtcvE5mqcXiollNpAnjqSl/sYgpRSnuNNkgFGdySWGfLT726mu1jL2hrdQswU2/q0Vx7I8
EnvHPf2bS5fjeB8u4wZULhhJrXzBDQATXlPpY43jGRM5CQIwHBfHvlQjm/vmDoI1RqWeC6dLMDUJ
3ZUcZ2p8L8wToKXAB/GeKo1P8KN5RcQDmYYfbMveq/vcEchEIlmxRC9t7u1Wzr/eE1sMn+Mu9jvC
Molw4DWKSi2Tlgk94Z4v+UEz+hT6ibtukXy5uYhRzhqXVo5Jf9tvUtQ55E5/CDWEH+Bs3bR3BC/H
uYvt53qXGLujsHpUaxPN+sV7FmGT/GriQAdac9nS4GJkn8gu/h9Zc4Z1jTl3Qq66vwRp++YoghFm
v9rG3Ur2aTWCodCZSG4iehCRaQjwTmzYJd387fi/tk/MZE6f3Cm9uHP1+4KoYj2iOTgoi5eLOXI/
RGFR0KATKK45IZsyr3BtQEBcz1EipLDwMOzvwwFh5qQlShVDPvkQ4ugqpuih4zIdTW+AQPePDc7X
qyzRIjHNwc4X3Sd0tT8Hxr88S+6P8LqLX0LkwR8/dFIbzVCEKaiRSn+szXtQp+wxx8J+1eErakeY
5zr89y1gN5y/l5129pgEiQFNBaqzWhpjYQ8I+LaILEuUyQWDnMwE2kNt6ltHlsw9BhSdzshq80Zw
TQHfdaurhyifqPRKRP/pEhUOvnMOUDyUs20ZYVmWIzfU/OPk9+nssjCMf7R5ZSF4WSUOzOrfwW4E
dfKvs55cmFvKL2lQadjrCfrLsUiq0Z2VjJ7QUCT8nCDOTMTjlTqv0pclBQaxrHT67LAt6lf6uKtk
G+kiolK9hZ3kSuD9Pk0L/06W3Mi53M+53V8meIV0VYdr135ZJ1neEJYsPfWTkZz/BLAJHPLN4YQM
ueMpka63jV6aonkL49h1fIxDDo+My/jwFRv8o9SDyFDZT1Na52stIPZX+G8DzFItylDdsCO2QyBy
5qCeMOyOWbvmGS11I+/GFTCH3Xlj1R2pqx9r52nPIhv6AD8FxI1pZUl2hPPl/Tsht0dCnNgGdJ8j
M5SCjOeK1Kk9htP5hRcsWgnPjQqBNr+0/aJouD3tClV9rj1fK9JVwPMoNwCArQ/SPaWeit4OXE0e
CJqEB58DamDM4MgckaGE9134wC0HND0LPUQWS5N1NcEQNTXkwbmKKkxQl7siqnltbgRTQLbLTkTW
oYrOe07/zPLXnnJCq5kbI44VA5oDYdUAgE9MwqFrnCFew3O3IospS7LRXrmr2k3BpxqFdHzUmJ2o
lqH+H2uYlu7fjEePVWYwFJt89SEnJpay0Fyb48UpA265uQlWMAQxr6qSjUicD2mDbjBx3prtHhFV
Ka+k2Vt4CmbmZcVv6YCe/UqxU0nB2Pi/I3Xg6vReOLqCZOCyPn98MCghWa4aYm3OwU0fx+PQ7zss
T3vaSQx6KsJD6K3FXk/YfwQxlZwrZKa1aw7+M1D1MkQTEcDp0WgT46k2e7cptc0DbWtRB6Ya7LyY
wrPVlr5AlAm5DgEL4iLEMv9fAp+XJepVZp/BbgJ0ZFHHJdMn6M6w+XCL+hPyi+cvp255QMnI9gEm
W6nvyeZ6JwQvozIoKNXKlkbLjCS9tBZbXKUlO8roeVb0dlZ9UjnhRNRJZ5srkvZWqou9IpE9WGQz
Oqx7YfiABLlr7yribVa/OhSnnBv+Mt8dHZlntzPDbeei1Sx8Rcz6P4hLT3aORbmXF0qVWGHIe5p1
iXay6hGst22lcIBjGn54B0vwjt+yWObRbGmRQeEzsO8rq7urFbjekWwg2zKlTxXq7A7F91CnVilC
Hw7tniE5N5rIqOLRYPLp+O/HvsznGZeKlrPP7/LfiErIHC3KHZPxeGQJOAQUDok5NvvmVOIGBchH
frLPBjkTRsSXp6fYYqVAkoLNCbrzCgPswnII5CrTi4vcRyaZQppLE1uHIntUZQl5pDIdKfAsOJCn
3NerajxSDke9jNEnPUD7iN5FiCp6K+gZxTvSDAD+ZEACtGmplh18qNY00OWgNJ9iiXQ63s/z90Fk
udfKJyan2OoQoaMHx0bEa0WCYp5hLUUnLnDcukffUytQ9dwjbGmEVqHzSpKsWFZENbq70+grmhYK
6WM29q1paXfgsMr8AOgiYJj4xrE4eFzKBNik48T5XQaDz+t8RFOiquoynlA9L/zmpcG5Vf9VmYfH
w/PzY69RewTOm2tHe636lLu5NrTO+V46HrZ/fd66m5WrUlHQc3OyxqCPpKiGm8n17YIxK0R/1H+1
L3wkZcG7mlz4AjAmBB9mqnTbVvD/pJig9770nubTS8h1SU+pV1IGPHJ6Ng9PqhbwSbcpw3Vh6jHk
OQd7CPT+VgWJanNU/4jbGVVxB1Zu8Gd/ykoQW/Nvgcilr53IXxD/V8nhBlZg4B34IdutNDjyLlEK
CPigoxT/e0ZOJfjl8OMP7xZKrLAQSDxfOo7wkEXlB0ZuVCB40zY8CyadiiNAHbxj+M+1FA76VofF
yup3DjHQh/xZkvs7/bjiDOWxieT1kIzPsdGWlro7WZh4x+Dr7fRDZh6wM/s6lnTjo716Y7/iv3/g
kLBozsNT+DYKYjMTzX42VW18QYd4fP/z1PKZKgQKrw8P+S2eo1hQ6M/CX76Pmx9YMX1w4q0D8cCZ
75WlgK2VV9AJHnqhApjx+SgcfZAACVFt/y8ShG4HEtwCKaZLCjVrNEBQ/LUctpvqTdkDtIIQU21J
8uIoXFw1SbKn+tLRwAe2UOZ3HO0kl2doMIfwtPf/io/OCQ3huCMmwMLgEG12xfJe5LhsYwAiFEaM
J9fkf8mTG88qzOFY3YWB9QOBoRc1eQxWkcbxFe14rq3/mzFEv69VQeb5ZgbiLDFMrvIOIjrLEtjj
f2a+BF5Hm/c3soRl1K4+Knzj4EszElQn7Qx9fcQpoZyaY6kfUzlH6BRKd0zqxhH5UXXHms2c7PhH
9KCI5wL27zM65UzLXpXd3qx2WAsNT5Z0RjLoLaFJMMpdMt+MTZRt9eyD38unvpI8VtUmo1DEbgeP
WB1wgzvPma/WSmnBQK61C6JS7s3Xu7tryDamaeCRHZaq0btiOm8pxdTNZ6FydF0euYgpnJWZ9myC
YLJy7b/O3zu/2JJUc1Be1IxiRHEYkSXU/PFKWlL06rtOPVlkYoHO+bg8AVsd7qRvAPO8KM0pqjy1
VcKxLlouMos56KQowOeBAWlVTVY3CYoK1moKM3909ru7wpc8VIPtd13W/XgBaUEKTJjnnZ/1XNuN
95a1LB1aQI+ZRdRGJop71O/EaPSH867wu33Jb4cBzxTQDcKSUtP/JZTZaS8PWuZV91un692BPnr6
b9Bz3B6yHq1rEzLL9rCISmHMnIRzUvX5Z5TZjyi7Jdg29J5Vbc+I5bX8OMnnU1VdRlVcqko4H/Qj
kQi7XXqXKZZF12ftoKJAmYNfFB45Yf4tzt7L+ryy3N9iA4wFzpnTRdGkgpBZZYVpjz3VD0zXTR89
Kux9HiRhDbR17DVnGPhanrnUOX7J/y5RXvPYVD5jMBzwuEMfx66yF597etqi2FR5OfsY4omLVMRn
wn0cmqfgo5dhIAhkqHbDGRiT+RdZ4+a9jUtXO78qijcOFVwEMa94Ez5b95XmEfd6O5ppULOoQmkv
YuHt6DmG4iBhYwH7OtT2ff3SSl1Z0zHGg5bavz/1YXwTIUbYsSHKmDaPoW0gn32zGy6J+F5j8K+N
Sq9CtXnSA0akwZlzNiO8FBBI9w4QhZnnQNNXBdjG30hudnLmF5EgIRlycGlgVN3H3dc0rMjLlNeB
f5yzeGZHMl+vL8//eLIoQZd7jr5ZWLvKkUGDYaXBHCmQnfKuNOaN0tNdGYLAWxXiM9qD+hF0+bCs
/tBZQUcFE6JoeUobEWXJX5gqXcTkdzjWbzvIA/0NQWx6teF7VSO6DqyYfSbOh5B8P2panEppjvSs
Fd43pupgTcSE9KOaTbo/GJGMqfVgR8H/Z+RWMurcEWevq8RTvWSunbhjhASD0uyOM4cUIwTwi85H
bzTRytjNGwocTQucv//wIsC9KORljAl7+o5l/il0MzWIgPxbPSpb3fnD4laohnnmJTbv1u57wPrv
h58ppyqccFG1n1SIqqOGgZR7wnczAVd1nihhSP81OmOQsr26PJxJeBIqBfYDlM/lYZZEePO3fthq
u5bZdT2sugAgYMXySDnwU6A7dkKSbvuUo03fO3/Xe/fKitGsLAtDhsq6LFt2EIim4oTetj35qWTF
H5p1OVDubZdp8xCHJWankltK8huhxBUwgKpX5bqXs+hJ7v3/S6aVh0v46axCbJ0MmOPPgVfRw0vJ
tuCCsx3hBamvT4eXheA9OuJ6HKXWXWT6dkllPFRKOay05T54RZbfnDhiz2Oc/RbP5RFxRiMzHMOp
gDJq6kYr7yFkGaVVY0vLAzM5w3G0D730bFEhY+Dk3Inp4CH1IFW1fE2kxu/9g3feWyCSibxBX49F
Iu2LyN9yRoEhxtIpCRimfpWQLk8jc7JjeSiYwHyTnarggvtPtf+ipDiShisr6UihOexlVxf2iFsv
44YG/AE5pknF4miZtSSwpPrjA2g2yOHMlh0Eioy9Fu5yvlJKGGYejZKe41gTdg6DOdiPCPm836CP
Z3jeQCsU7lWvfZV5RA+JB3b9Q7HUe2CmfNjYquwKbn0xxgNRoXHbAO6n9R5Gfo5O+rlPqPlZL5dC
ZwDLLJQ7ZFfWZHakITsMFoODaRm0iO5jCOvwEmTf6sXDuK3gRyywlHflZ8yYkSIuCwRXlZYMhHEt
Fh6W7AX02Kb/8bOnhGhCmXF7mcnoj+eA4vrJDGVEErS767M1A5V9ar4vYoK3CNknuIC61Qqvrx3f
pkvpC5L4VMEHmvPEyKkRa7sSi6kGqCvyIvkDPM6fW/kpuzRryqA+qmtlEZbanTRawnjR/6HFmM5U
kDKOXcrGd7kdqIpDCSSZ8XNAWa9207PWSFDLC+zGxCssMaJ6VdVgowNL2dc+2MCMF+7OrI8G13we
wWi+sgHmgTAclWK3OTFkitDeIOUs9Zvbabc6EpDOZoy5CFt8KoBmG3Lz3iTz/6Vt8TnPn7NKcA35
c+Ig4v8Q3HJjMTWk47ZrX5z6xK78/flazR7l3m2LVw0zRB9GULGloyMRWumrebANtcpded+S4fch
MY2i+Dvo4e6c3Sda4S5gyCXCE+Uy33QNSwKhqVR83xyIfFVpclTul6dCnAgSJCDaRkztO+aoI1o+
1KhayeNfuuWTkGXlxXjgy+mWf5ah5MYv91+k2d0j/6N8/Pq7+4G9WQCmTe/n/cNMn7plO7f5HYkV
3oJJ8HTYqZP5qY0gCQh51jjzvYRA7+m00a2dwKwfmnvN01JVlZiS4vLJgkqwZUeSm/w27jdZ8YPQ
sEWZRjHXPaTL+PF5PydFAyREnpZnCxT1OpcsU1Vydm+z2iTshBaXatHQh+cjTPIgRBFfVzvfHRG9
3PtA9xt6X+Z/JmfwdXmxcxMxLAE31i7V42HUkohobXQnaRJ8fDDjPsu0Srw5GtzRucN9j0xzBTC5
zy0DA8wWRwMW5N0EPrei2Mfl3eSw4MvMt3Gx2dACyLLJ4tAE/XtIg93FjiAHJoD4zsRPmjCgsJ5I
xrGugd8ZjZaS581oM5IcN91tgCAna+1uDv7OJG1IMn0JvZ05GbEgPxr0+dW8srk+6pZtphRfk0bD
zBqi9xp2hpT2qSCMCy30Ld5hq83Db0On1+YKbSppPTuMz2dBuhuYOgOtjQYuq6PFtyf8ZWoJH5CY
X3ZapfbWgvEPQMobSvyaGnKiD5kq7ll8WiXW5FdBzX4Ch2mPZUp1E8vpaIlpFFPtwuP6T4g4c/h7
C2JOuxAv226QrJbsG6HO6x9/j7Dxn6gD40ZXHuACkIEzK8UylVtz665LnLWRyrjO47DOK5U4kwws
sXZ/KZMaTMvEe41B6elGY09ktrmIBt60apFXYQeJHxE3Zy5OVDxJWTb8env0vToL5k3Ls7ilc2Oi
WKBLmhZLiXtFUPK9ZgUPXyHqM7ykSG+PD3QKOmaUSDrKKyefMzxAmdFQPiop0fTF337ecb5Oc8GA
+KTC79pZysWOFijvX1It0xWf9/vzKrRwifQWGr89zAq3PiSHM3/LjuuBGLf2w2H2hCr+9iwbUW8P
2rgq/PI0kFwxgyyL9pjammP1frcnIFdRwZORPkC8nVDdGTbdAnbMAhbLOFwhRt+7TAQ72sPnJFj2
IUiKLTsdykBbNM/BniWjWu+Vc7+nY/QgKPZUFasZlkIyC0jXkG0xxalbZitXYCrdPQvg6wNcc2P0
jF6a8f02hLbbJFN36zi1eefvsrH43AROKWI+8C6PxNGug2vxD5uF07KE63kDP1lKYFOaEgqPBS9X
s/A9WEkYRXZka3knqu71S80GPp0Pw0A/RawPEJF0hfokNi8PEhvIqoGkfSxB2Hem9kIxRvWpoUfk
kCDCPjxl9GkqBIn9xs95FfUsyowUJ7tIXMUWCi3iHOtCqgEQ7T2xt0hVSYWF5v1C1N1jzIm98u4x
0XWIY0PvLCJfnyFOSN4Mv2FS+zLaaX/u3w7/oIJBAhYYB4UfBIMd7p7+XgVoVRBX80CrQbrFcL5h
0KKk+JxdVomOzqq0gX8iS1NiUGsEByFFvgFCR4dAHY0j+c1Cw7Tux5KFKFiDw+cQAHLdmZ4lzwDA
OMc0r7UTCA6pRDTcOo2QkAJFmO5qZ+j2hVJSG5T2L9v6kmUUIAEE2MmEfw7GGrX+L+CdEv4CyIyB
MOcYIYcT2al0XtboTjVAOKLukdyi8o1V2bR6cTN1BCL6ubaeffAut7PuuZAUnn2zrbC0cGzbGg/e
O0hWcqVyN2jEjTNrKEiGhRq3GTVfp+T1wB3MsEdfvCpf1fyzdwl1KbjMHzubotVgjb/Uh69oForJ
dd+i2nguXLx0DZWX3AiBhrZCUjkGMCO+I7yCJswA3YfuXgIOdOkf7Cm5j9ysR5qExm9mTZw+smxP
qmjZ2rHRaAQkBCIzKhSSixFD6XLmTzFKMf0S9fIMvtuJ+jyxpYbJEb74CTBJaQ4luVN+AdUHwpAr
/SgtpkmYHXKzb66JBsWqQPUjQfKsVcw8TzoWOVZpwpdeKRaBJSQoX+PC+0uR4ndz9XOsZv2ug9Vx
mO/fGvIVAolGMBN59ifn5D4FAW00G7OaQAEW2a7eJDvBYhwkbGchHwCUOlyAKDQUGzkqpsaj5z90
fK+lxvo8YF2T3JMRK2uoXqc/0j6Dhn/E5H6a4Ikz6nZf/6Z1s2YT7+yhqDF0my+bLKgjozPHB0pg
81PcmGrDQSEymt1qE7l5ZpGU9dhgEtbFezLm6lodP88mZDWixwC3HJ7rpzk+3lEisUH4+8hCOE1m
3f0Bj/Wu6jmKesQm8/asiEH3G7F8ctlH8qsMFZu/1KUDKJdcB5GCidaSRNKHf2QNikxOrkmadKF+
PL7vTVuhtV8HkCaZaZ+ctzDTdK0xxfftUDKJA0kUD+HwxRDwDVLuu3rR1t7CUzBvULEsmxu9NWds
rm+Ws3oGVfw34n6H9joYGsFTW8BoF9yaZdvj1xxU5/N6aQtHWu7ODtDz2O3P+WRZVb+WIhxVOSHJ
L3hgBaYPax95Yt80GtQwQ3yQo4ZcHskJJOEhSHl3dKrFuaWDhk8p5L3165wuAG4SpUQ8BdEI4e5U
SN2mufagyUORI+Kgdw2vkpHoIFItEvTHldby9wiiauETS1dygDW9UG6G+eKEbFQHXIaT1FR9B8NO
Px1gPfqXrq+fve2GE1S8PnTJpW3e4jOagyGEZGUL7WUoSSjZXeXxrxM/joY371BT7P2azVhgE+j7
EqHrmasEP0AwTcOCaPUN6P9tzHvGnSu8Yc9mrY4bkR1kddeYE1WpJbI+GPERuyM6RKe5IxZjImWI
r31PRwSy34dT46SQ/rj12TOOhsJYxTnGGaPPfTwo9k0Tft5YA/BmQWIUUSolh7YcOe7bu4WkNCeI
ElrBpRzAHqOoisGjbnbvkPvcn9VQfipMlhQtA4qzR+/NwSnWcZVqC40R5DnN0rXHzu1c1340+6qF
G/QvayWXSSyFhIlbK4RxI1Y/BMn7IRUpmLsI6hdQZPI3ALjzWq6FJUArePJPTvYD2ljbWnVzwyVo
YvUPAKIiT5WX/0+8f/M/06Ed5gYK+bdq9uZN5JcX3iB4UT0jeczLdODfxaj3w5S/AukK7+ZF4K04
j3bVNEU6d4z6Q4WFvdVOmL2yE2WUe1iDk/QUZ5+yC2ENMh7v0kfbirmmMpL0ECk/nWUNUqnOnvxj
O3WxFEkvsjelt9T0wXxUWyWD28WNb4ROEsm/gOOJ1I3a3/o4sxV/tCGGT7jUOGF+nsCMEbn5i+uz
N7dPrTlteKhcSJof2aEU9FD5CMMc2VJ5B6W51G6h5PkR0QMMB7p5cbb0Qca4YWWBJzGp69hjVpq3
P22R3iLjVmlDLCz+weO/Y/MxkZqmqq0othHkhBayGDsPBiZCSyyvecacWj8l7w2aDW7DnElnj8uj
UK0ojft9DPsWo/6Fo52vXwD5CxVzWCfZALlRqDf3MdDU2+jOUucYS4ehBzAXU1pNtMJyW0vy/2y7
NJtc98CvlKE1dTbjVN8OaOicdgFAYqsU93Skus1R7JX/zjzF29xej/8sIo7pD/J2UntJlAOYkcZP
3rL7wJDI3wW5xPCZYw+a/St4jAfg/OgggZ3ieU0Mk4fqo5oPSa7HLrOjF4zbH86EF6KqE2f8/gYx
S0suL0+tB8esulF4olVlmtUdL/8NreN9drdv12/7CWMhfiWOZ9F039GnrZru90bS6FwRrTsDXTuy
7ZzJ3/FVWhh2DQ/N7lpiMvbencrANzjBn3y3wDHFN2FDqPfp+LqgL/HE197QE/5MNy43SnErpnMb
MVSZ/IpKHokvML9vdZLXZVsa3j1BZodMmPesLNEr3E2iQLsT86k1U09/g7S2R0RU9UAheW2eBCbc
gexuB77e0cOg4iagB170//5FE0FFiV8rokVWcIw1pqizKk1RtpFRxdBYSLXi9F8e3XuVsEzXgHtM
zsza7Ue5ZUs9fwDxzgD4ivKn3oOEcZaj34jzC/u02o0ownu9yYI+0nwsIUGguksy5LuvOFInVZ5A
kiUopOBzqbwtLAw4fdB04/ARDuTw1Ziu12zUTpLR9PsCYm5UbBqAQgD3Bi0WL3ABIEIi/OFmoWNY
T6tQeM7u4yFEf0J0nFNuKO5a6R2QmuTlh1v0eb8VEp9OvmYK8j4+GolvXrYK/+wiJqTugMT0XgoR
ParCev/LPd5n/aNjGiCK3Z1dohL9MRDM03vJd74O1FFxoveICvlFlRkFuFqdg2vKVYgHlRdY38L4
MoXVNz2rEP13XRHKMbCoobieB8JnWasdXXkshb5nXJvQddtnnZrIxNr57vEdq8XGmDcazJxkYtDG
Fyvt7xACV1/ix+SCW7WePp85gkv52qeIHmaXXp1hgP4zu4pCMD6TX9TARzu9c28ynXRiaBmqGC+n
Ntkuql67eAM+Ne3LFngt+q3XOFpD/1n1O6zl+ifTThQrtGchO0T21PauYzm1n1Hv5M9XQu4Q+yLd
bOk9dil7C5sGQ5X8W2+GELD2h3XkzYAH69paEs0FptPlQZIgh95UxQkUREnAOHivWo4aM2OFvOqL
IdXVbuICkc9DKivwMSYENtAPUH2A8CWyI5WuFoWRYy+VjL6kYTiHy/Vg6w0WjJ5+kYChqzaj/s1z
5mxmdxx+Xh6jIy5A4cnUVQ8t9rE3R6eyDC1VBNqOhAcLRAe2R7MgNEypr6/Wi5o/7UHiCuzuh7/H
kcX1uyfezonG6uFscF2UzmDsI5iJrg2+cHbWsQOD9AUFuYzXwpd++qpDHeVOC7N0PxyHTId7kI4o
DYJ+rOWZt3AQppyEwYR6SfeWCsTIdqCps/Q4EEJyWzJqzYWzq//XNQ5BTf+U+o90nM7dwEACaDhT
vDYnxs7ejAWUcHTcrFLGBeJhslMVMbwhN5mD6/qWmj8YvEO9SFGDykhwmvvCBUPtSHIiUM7pL0Oz
iXsDVAJxmZd0V7/TeovOi2j3J/tJh7WMUbMIA5wxGda6Y59P1RtsN+GNc7m7K9w3BQpYjaRRwNgg
4EjMmdagugoQZggTxG8tY9lIga+yQhiAn7e+H3OgE5Sg6Qzj/ytIayHb/0KGhgWq7aj88HKj4EG3
+91Qd1pPwX8aFRppMF3ksnRiqlsPFyyoVxdImVSk22L5nkFS/OKMWi6KQDQruk13LlgL9MyU4wF+
46iBu6Y+W/DHEncBX3aRC97rSygHKCv2TnQKFjKkDbzwUeA9I7O2GfMkTk8I4x5/nQdtAuzXADdY
MVsAlRJLPfDzj5x/w/n1tPD1G3RcO1TCnz6Uq7h/c88ywm6zI7BvbGgbMhChZMbwsdFIBsWpu9LZ
9Kej8k1t96tj4tGfV3JlCTRbokTMmu3l63dxyjmWnALDAd5QD3ADy1J+Aq2oZaMFFkZ5EqM3STKe
yFhHsHNIP3WDtR93NJObEbRpU6VR7PqY8UQN6LlE2iXksuou0TppE3PmssZtODt7HqqskC4w2f3E
LSZnO1ZuPefQSWVyPT1h/YR97w0LWaCfWqOdxYFfFysJiMWXzLo99S0cmJZtkcFhs2GeR6Dbh8GV
y+dmD0wMCTQVGfx0xjGURZ12HyrSCCCGhtEXTWgk8iJzk0vh6lg1h5bl+eHclqqGjHbQoUH7i3ZI
WmfkquTOgsUatZvzCNyHGPqCya5Si16Gw6p2lG6BivKj9pItPvO4enbzu5aD8GkMEoWX+wCm/8vL
uPbW4RqAQD0TtwJtnpib9lrny4hg9BrBwfUQiZiV+N6D+bK+1oglx7buJOXvUQ3NrmoYuWNra6Kw
RQPULX4aRbyoUyEwsdJshsbT2tczlp1UCF8gEflCKXFF91purn5mqi6ZrMz/lDAlfb1joUVeApHM
ynT3HF5E0brFsrirFxg9NlYTzSukQTCU3hNA8iTE/5bBvaaeTRmia9DW+dHBcR3IFj/i2wrsC0kr
yaCshjA1byVIKwf/iraYg2dibXITK+ok4mbi0cZRNXbwAZ+Db18OaStOUR431eXvIhOTaMgMXoQd
j+EyiJgM8qk8R+NqiCfw4t+eZELcQb33bw3xuXwjXnDvTd9aKSZ3DeV9leKrpQqgkMnGH+lCTx05
lpDeTkvDx2JZgLrHCcwo4xiFyop9Q9eh6gCNIbNsVwG4TlsLevpq/FWCGxjdJ2c0RZeLLY1M1TxB
Mw1sF4MyweiZIXY7WX+UQNMBLDOITtyXMWh7cISjkqdtmGY09FLXGqrd1AFbBN61ItXkaP0SRJL3
EwpaxUHgAGjAbRG5kZDpAGYNzWGf72BtwRr5jllyZFShwoyljs6Fh8FFjN2DgsskowZbATivDRir
XV52xmkYB61W7uTlbeNsIzsz3ZdCAsu+BA1EYeIROPhFvEiC1Zlc2bsX3u1BjSYN12sR31OmujWJ
AOwV1XqXPRwMY8WvKukC0W4SEcox684CSOrWxu0rKvhLhLiNSuJ0bfgInPnHD4M/CWMXW1R0kI1g
lZ/bs45SCEXBlc5dCNALIzGnTGmDFznBCT1avJAnL7OJjNHqsXv69iedgXJHurxTTm422stRjovh
HPdeNDW0p8ur9nCgIHIO9RFhtnMDkT/LPFDr7b6w+gv8AnWMJYeZVOvViuNhM/r/Lkxgiuv7Fs7i
OBTQAKNBaCVKrsj20Hr2Xah256zZFW3b+di17g1WIrwOziiJJD5x3icwn37bUS5VVQnkNsL88EnR
GBx1AYojPXlzRQEPU9Ra4UDZLcgiHUsvYFzkRuXObp+wmer1U4hxCVtuh5vgUL6p41iII5C4hQ0n
vIQSPDVVlO2NXOVzJGpT0pobI0h94mtZdnRxTY4go1aAOElN1YvmOoOdNiiN1h7CyPjoXa3prTrQ
4unJe5jYUmX/FsEDqVCUvpphpt6yyj59fQZmjeuBejlx92N5GEpdgp/be3LevxiBEWSBuVVjyADi
xJwaLYET95HZKAXx8TXxXf2YWaJMutqs4jiUqL7OoY0f7zu9/MVfGQ8OaZPI3fqn/hnN8V9s9xES
UatsZNvoYeODXVd5HqazG3InVZx+FTPLIPO8jqlgBSlxLDjIH7qnz1rnnu75aIgHPTRfqfrl4B2g
OUc7LJ+NbqkrfDvHyNfH/uVWNEoY6/8g2Pwchfohil6ytSuzuKj0SKGpm8qjj0GSGft9pLWS3TLm
jjGsgjkmzu3m9THg1O4M8Rj2ws0YAJA38XnXIsM5NqfFOAHngdpvNphphrXnNrXgbHS2nn+bfYie
ddcbtU68t8ccDW0GsAVyGqgSpAsDA9mu2XHH5b8e16pju7ncFWUB3eWwolb6/WkFJRMnPo2qfPdH
MoeasJ0/eOkcs1dV/WaBiwoqHuOxulnVOWQE/cVEZUrJO3iQuO0rxHMjYd+SP7jCK7HjAJtPcAB3
YUDrk9ceh4YYyiFf98BZAsYSAIz18D3VkfidZZmym08IIxQ9FN8/ZpjrX4ltcGCEbgLHKl6EPLb8
S7UOjleb46CI6uPJcOns+Jg/fLlSE7ToCg1d9rAVAC9gmuApjOJJUAnFEcjcFQn+jgVRojZbxHwt
d+ERL++vo+NkrxJ8d1vkJTKM6uWS+RSa92hwRlYyBAqb9o4T1HPJ3yc6DOhkLLydzKJ8K2a00THd
B/9NYeZ1qqTXCYcTQrWltYubvZpUrwZlq2wVCLIwh0D4hpLfKxaZsj81RI0ImcMPSa6OSDVjPVge
GIwgWYqf3Ej252Vw/cNf6+W64Fbw80xIQiilwIm7aIq8bIJhG4Y1a47emCMpEq3/ThzzHfDNN4Vl
dTWVb23gzsbaCrYMWgwrneoEuk65EdldflEg8DdUg5e9IDirHlxDmdXdQOs5BSpxfDGdjBFrU/LI
XxEq2698Px4BXckTgAL/rnFLHKsLXGst1MZAXTUD3wPa3b5IMhgmeyqHF2ElznGrxBMY6WZPS/Fw
I+WBmHwRUDsxzakO+6N1HSRGu73NUUx2CbR7T62UVt6AcdfoxgiBitsbQyCpbZ+Hm/iFAey65t1H
quD3avRO4zSYnx+vtStLnQrWI5ceoeQcIxlmbQ0rAvosfTsMC7kRXBiutbqHxbc/S6/6GEbV/nPg
VuK4fFxlz5VYVSevQZnjZRnrwSZp7dglqPYZNPLxky3wQ2ohviAAFr0RaO0NvLAeDXPfGX7Uc6fg
QO+3rWdUIzkouDNz2Wleevf/bBeowPrV0dbz+bsOOcV1km2BpK+3TLjRk2zwZPWt2dw3wXiA4VD5
R9AlMiMhYc3EHb8tCVOVQM2qCTJDfHfQ+q2ufjsqxR8MrzmHAcC7cq/ZyavDjG9K32UjFM2GOmI4
ToEZrYsUX7WDNF3MT1CQo7JUqc6TRiGOlcYKGS/OobXvtUUYnJNX8qF0mYx1qU267oN4GG5whA0Z
1O6iZ6n4qJpTvTsiGxqohrKA2TSqJax6uY3tHDPAZn9cjfIc9cGxFNQLWHdEKiLnMSsAsAXa1QcE
fgikl6qUeVj5BbfThjzuCzK3rDm3UJ6v9Y5U/o61QR1qTdLhousFAhQEhz2wfSp7Shp0HaIPpcWu
LT3eHuLFJtacoU6z+pVs6UZnO/bOMyujyD1qHsmyPUwNQ8qROsOzoIycY7CJfybQsz3qlLV9AwMA
V21sR4x7u5WM4TjnXCktmvT1CwaKLPuWXxQ6rnMKwhKRw3gL+FKmSWyT7LdQM4PV3M9scfjFem7+
/pkSp2pahhN9liLdygo9q4UilxWJ7OeMIuTepJUXA7COpS6sEoCQqsFzDsPgiofNjCdADjOTHOeh
nDzhVQzYShhzCuXB8kJggPzsoXUM4ynAXSKSIPKZG6PeH5DGnpPSf6DUxd8WO0BVfk3LBWmZAE0O
UylUXREIAnVkenTTnZfyg8LZ65NogeltRam65JbdUcQXWFeRCYO4B5TbfuD2OMQtANbpOel9U1+7
ZFKtpoZq1OlCtE8Wc1NEbDt7EmTuvIMe8JRx+GETVCjGMBsXOUsqAhweoCaisUTuuNpWVIc46ft0
Z1Lv45KA7oxdZ1ubUZ8sTG1ZirjVzNmqICDDdpQq7IOVBPfPY4ZZmeXgNYLOIopaDla8VAJKAUwP
1BMDtVkLmZzfi7w5LNEviZYYfFq0zTbHbpA0bxBsblW7LmDbjBbWOx6H5uQvAu31oV1cumBkuvGi
06lviFbhfVKe0creicc5zAOYJKLMlvzYUogrcwfyCM/xTT+9zs8qzMGGJJu/hbcI9WBrqlETDzK6
0fI6b0H170EF7ViPhr9nzlizi/BJe5DLf61HC0FGtG8FaroMXSvZCxMytIoK2myHuvlT5J13DItJ
gcDuDZZaKxWbzr4P+AUvUSZG89E/vhdJ/wg252hU98XRWnnVRr8Pvoc85QvzIZYzYqNiX8WaPVik
MA297fn7cryoX0w0DtFIFF3/vmHESS2dvkWVGLP2LM4cEueQ+lt2St1FKMDHBMPhrz9nxe2HMde1
43tdTGOCRMUW5dOQH9+HHo6fYK4BZOvx10O5B7DDfhY8bEkotdok/NyDkBLxY3a4DSlxuuSi03l+
DhbhfkuPPhG2x2hECV95fjIumnlUDtUw1pK04Nn0kvtA5mrXpsShgEb1u+NVDtDFJzAvxm9GJL+b
Ti94JsCJWgJTVu9HA7lT7sy73//QbsbTyXCSJcsnWP9OO0BzTXpCAJyS1OUuHpTJiDVk28cfmONV
Z3Q0gBZ1fH4ss5hdL3+6tMkOLuQILB2dQRawHs81EbVsOPVwly0vCxZTJIkKT88vn0q3JcDmD5bS
GEbNl236EyVB++ZwlBd88tquNsJfUrWe3GsjcHWPyImNWwsjA7ufpn7RWKJviFUCTJtH6ayQthU0
bv6lPmDXflhtNbwUQK7Bh6FHSiRNv/V8jpeb7lJspu2qs0wt9hgwBc/JzD99v901JlIht6JcXTlh
gEOgbpvbyjnBNiJIhemplH4YeWgiSDgtxalh0wV6e88bWTDNnFJqPl5AoHf0WP95212Q/iCDxDJv
/vvHsfDiB2TBrbd5jZcNka9qKzU+u+Q/CB6rLU53VvB6rcrhp6YzdpOaabmVaIUo5Gf31/3XO7oT
DWTgRQqTK0oYwLfyzj2szCCgzwLW/YCJqh92HOOJx+kgENkML7B+PKD3HvJWpd/QtK1+zOvVmEX6
VUvpYCyNi3hLN1TgsGTGxTWF8Qs2jtmJ8AaZf2hXFKgwXvlUpMQBhmP0TcDkivsf8MrBhp4qPS3m
5A9HVxdqiNxAlqkYm/5+p0H2p8eAjIndKRHIGr3OtHUM675OqgJ6waksALL07hSVDidy2I1AQ0Nz
JUw3hbrB6KO6RqI90ZmKZAtKQoxLPg/l8XIuz2f1T9P3OxpM3vMkePF5TmABSuaPGCYbrtib8/Pn
nHCd+D8O9mx/W+L2PgVyPa1/AQqpXWt0NAmTNdeRpbV4bW1zRootsaE+hbarMM0HnjY3sn1w+JlB
0gEG6E4l3swREASpSVL3PckTwhtwV0xm8qWmym0Bj+57Dx8foGA42dzGz9ubnpN9j8GmuECULwJg
T8kt/6dyOIoRsogFPxLMP3mGWeJ0xCxLK1rHug9NK+1bK1RPOUpjl/Zz4elqrLzBME1awYXdZtrj
r+v2CIJTxT6qs1CWJjEk9G8fO/eJi6ElNkLw2dXamCgAe9RfInVAW75+fNaTvh0fquR5jEVpvdRg
Zg0cXjTgcajGoN8qhho1HEQLCvgGV8H9sV2YwMnCPZDSt/Y5tB9kRXyN9t+T0wFcVeAlaen4vw8j
o2FIZZ/VAw8rcm0+uDj28xvlXeAbH3y8/VCjxHlE7/z5aqERYmJPFs0tuThD9fH+T0zQBIAkgzxN
/8WcoQoUQ4ZAoMZP27li6x8UAMfv90n7AcWmPcJDPX0Dfu0DCS/DwAZATUy0xfjcvs+eAWh3JRI/
vlDTASWjaIXw4nUr/ZA8IIAFEpz45R84xNgPxIdyVnDY7UcavYTfZZpxglguPLyu9KlE4lR0qnQT
6mVuMucEWzGqjUf/SEY3jj2uVE40LiWGTMWiqk/0D7gxdxF4XU8F6sLqpWBLpr9NupLPFhswt+uU
KPyYLl0/caoSUxBYxyUQJ7PPQXhJao5kbbX2HmBYq77QsEtJG4rRB4Hpoxxa7hSAbUTb6vBlP1Tr
1MzeIj14px0cQeQv1RRxGuCG7cdB0N7AWQcu2pkmICa/74OZEZtgScJU6fjcc6mXGazN35EM30Si
e6KdCrVBjsdJdX3KnZCMpqgphlCSfXW/3hCKiT2OADcae9oDxUpg6HRuN3gZic0Ji1xs/7q6p+MX
ypMXxGMm7hEQ/1s2b2l9ztr/Gu9vttgjG2vNa2tfEISq99HNgJtzNyEdysbHzkcqP9760LjoC8Dr
Fw2rwHUqwloH0rruWvzNSPGWLWdSE2haIAwBnfOd5cBNoOYTfZMMZ9GZ3q+DpJZwtKUvjXW3PgR7
4dS3ptV+FIkmdSTWwfi/IGdFosFUNQnUUcqh+D5OTBKI4iBNsfzvySDx0LOjfDJc1djvO6YblBVF
pTmtuNypc2QPg8HS+bzieotDti06nEKoYGGAFP4KNHQGv8QBnC8Z9m7JYZ2rAn+wI2iJgmT3LCct
9+/drrk4kqMGckm4zMbvabOYy5S7vF0WiP6fVja+LPcuennlJ69WC978CSf5crtDT0UqG7hoVL+C
gwiUy3ofPlX7zqMubxtjs4IhtihjNjLi68qwafZwImMHMYZJti2XmWEJ3fxbjTN/JkkAUWbH8jp2
NvkO265Bwyn7iSdk/SHV5GlJlTDdQkBC6W5h9F4hFvbNNT/RezA82y9ccTnP+dCmC8QlbQLfJHFC
hxWc3NWTCyIhGMQjVFCQ3kOJPjRBOYvBapL+sthCdim72dLf5DF48xAOApIeKULMhoG2fLSZKKIJ
b3ZJS/78s0UKr/mge39+6rhATCwfMirRQ63btZifC6I+phLPQBpP+K0NsjslZ2pz1HsoGynFIgHK
t+yyjIB5bWyVKorhvrIqCQfh2oVt/HEFywowUQH3yw2K1EpJBpU6w3YDTSFKYNy1rAZKYCBMCNOw
MYL1gzVd8KBFWz4JUH1e599xnj0duK1tToDXJ3riK17PLAEy6Jzep7kWaQP7whPEB53p7//HBC0s
2p/RWtuLWqVTNbZERN2yjpV6EOTe5yuN4bxroPPrvZE3WsR1fggWSp7sqhU9FOnVmuBR4zfCfiKc
1RUB54PBS9/rpAFKwqqb3+HOSNlr+n/jEzX/jSV0vsRLswCp0tBg0btIjuGy1Lccn+qjQCe8HAtP
Nscu34xJfqLP4MyzOGyq7xJWtYwhUp5CBmNVxo2XbDxnfnUgHDhImebJbGkV7/nRw1RjO5Ylx7Od
3vRxGrZB6VSQvafy05E5Ghs5RqUKNs5YbQWQvQIN7g5OfUPPYy/gpL0LdhgTEeYV2p09c6KLCWlE
aNfzSzIghAw/WhR6TCLdrRnJUMMRWF316+aiRkOa09Ljm1snY2GaLnXj5eFppKDRPQP+JHD9HCjc
y6AX0qplUFg1JZ+MonV/2R2j5quEUAMuIT+KbazCwjFkdWBWB4P3tLLucVDj49Ow3UohPeYRlMn4
pfzS6UPLrArIbgg6Lrg84IhwzCLpRIdzrro0CHHt/GwHhZFZ35spL9PDTlDuJeYVVxSfnFdBsAnD
G+xZK9v72sMoKaPSU0GHJRz90qKsu5G66aNuOawFthvw7ccgXX6Yg2GFBoqZ4mfjUyPJUSaFp2AS
y7eDylkVRPc5qqc5IIiQ4lQcy5IfzpkI78wWcozcpEgbxpb1XMccfMDAvNCzEZdnhA67DHTohChG
FP5qvVve3xJ+bR/oQG2g4qY9zcvRi9Gjfk97P/p7g2V3HGuidOeu4E/DMnxUO1fVoILUunnd55Cw
CkYmUFto3z8g94Y0BSmYyFDpz5+vo+IfTzH6k+ONVPo0oNjmODVfzw+GhUG/sKMZsDpTBeNCaoFU
7KkPBV8zaPcpKTULalRJMh+7Qi1lsBdMKLJufJ7RkIDvFZ/9wfc47ExSOpYYlZ5fETrYhQM6GuJV
zo7e5IbUOEtuD770pcIX7dEKqgowrQ3x86wmqx0tMi1Sjz8UVBpXZsky9DQ4fUrFICxSZybVlySC
wUGtmkKCXkbbyuG6B0lHC4NYrhVm0wZChwE++LfsZszRlavQ6bTYs+0spYOWoP6Hoohun+dZQsZ7
9mDvlNidXf6MEY04R11VXK25Zb+k9ZY7eBAJ967X2HyHfcIbEaxKCtSgtyicdkGVmUHDL/duKAgE
LwBW5iNqXWgpTzdyrkxTEN/XWwgKOppTAxVzp82dozvEHcjcfn9dEpu7eXtsyOW85eWcSbx4CNg7
mgt+eUyhlob8zEkzj83UeWEqJK8KWhvVvVcgD+Ew0K4zXp0vQlyBnt8aI820HldCg/eKoz9+3vtr
Z+zfCa1eUk5nH4Wipk54B8bczsFMF3SPrZ0sbbIZeexpcUglkO7NrlsGcuLGEtf9+Hl+K3XsQb75
vFD57abUc81Lrv/6+B8uzEuFZ50qur23ZnFQuXrtft/D9J9R1fwSgHmdhyciNVXQqTLwi4CapTeb
6W/hEecPhtZ0wWkWeJN7mVGtYaY7olOuvGaNH7s5dcjdqHG2nxoZFPJ/XGAoDR7WGhCTK2m3AtWv
gEr3coNs9VX1baTYxrmepCBPR9EdOInfmvffUKAzhi1pj3ub0rrmFiVrNBY40V8bVQQDxWrx9mG4
jj1eqvpHWPLrPnnjtt5EHRUKQKPt/RKzECZxYsc8svONZRV2B7YWlguV3bkZhxE4jNX8D3Rz3vQQ
7FJ1udeYgKtAUS0YP0Zjc9F9ZM7HHuLS8VU7cps9SbaYm+oj+6c4fzqwfdXpKc9Iif1vJpJODwnq
M/4gXoopaFmSqc4UU1HhDdH37QyMwhZFnHLICey0yAYSGfStTKkG6RLxF5eYC6P4cerFp0N3bx4E
JgoLgcbSnxMZr07azXmKxEnU7FvszhBA2S9MXk0NVB6gXS64KMM9gcOrJgwaVxyHzMevN8qikIUK
G0F+/sHoEm9M7KJwd6vwxMowzSvullWaSNXSJwN1v3DzUsP5/poYJiuJJMjvFAIlV92i4EHGsbvx
g/bYKAg/S1K9oQn//5xN9JgfqnBiagpYDUmHM9Ikz9COLw2ulYL6PIaHihKvlZYRgr90fETT5Dq4
AY0mhqqbbQF+TcuAj0/BYg60kANwur+MWMIu/ecEfuTYYn8XFaNslrMPdHZLILzO/y8wymj7QqPe
4+3Ny6GEi+wKd58gId1TjdLrVHg1qKotbGqClUukudJu9277jefDGkKURzDDussrMd6ksXgxcafK
RnGyU/jLpu0ngMiT3W+Ocb6UFDS1DFDZfF1bgV0904YlQhhko1c1F3JR8oC2gaxsk8fSL2TcdPnV
rL+swE7O4NbWM3Hoj/2W9ZNSnR0WQ2sN6eWSBOTyg1bMQ7WgGRv2iUZBMG5acnPWnQFUE7gzi/5p
JUs7VymcXruiuibieN0anqj98uQFVHte/axhR3JxbOljj0p86s7RFn14W1dChH3lmTJFqIddfoNA
o3nUuKVAtwZC8i0YA/I4s3XIRTN7RMwlxHkIgb1+VWAcXPUPkc8t1ZI0sdspTc/MUBUUdIaNrJFb
G1BU1oTZEVOuo73fkkGf0N3dbxYON4VcxmgMdz/ZNcUZ1EeQpT2mRt8z3/np6IJW22uZ8V7sKs3q
lc1ZWkn9eOgDNmRy+0OffZaL33H9AslOaMjGXfajKAeXzBjw88WIQt1KpoOFgV0XB3A+FjsmbK1O
sZ4pu4BCodhe7gyrPivBr1+cxO4g83yN4PiPjsOZgaN8gxDqajaCvHHcloQxNcl+fQgsQSCAibu9
StZocH5b5QFje3MAn59w5zAkR9yYNpPtZDQ2xzfDjTe5jfStsPRu29isQR+OuslGbnGhp1Zb7Bh0
dMFTXchRRtyF7FHgcasu1oRPf5h0psWHGx/sp4rMDDGVrkJgx8PX4nKaBKiMaQLeM9I0ohe0Ridg
44+QDnkHMJA8PLH2bEZEVLpVo/YfIzeAaKm2U6YOjw1AUwnLrW0er4Fcj/t76KF2cvewgaUNmRFL
nHFJ52kmdQiPyJlkVdUUxACIXi65A8e3pvIm67sUM2rhcLFJSYXaAOOM/rne0Fyn1IZ2cHipqInx
GrmisEAVgS9Xe1h4oq6Eudglx0YDDnwxvlROK44hpMFJh+aTRn2AE6UBiEGMOUorQl5ZfSYoWrUF
rMWBBbxaiX5MZGD6IwyaNJhDJXHuktxr8E39FKFON9qA0qkkeh88Bpmj2YCWrwKLxLcSGDRVnEO6
8BVxVyuPfQlXd+Emrj3+4CW1hT1xhiuBrhJxd+JP8YA03fnu0VYBRZOgWdHF8gnfSdqORjin1kvz
/ckw9aOez6NREtvgsU68Zl5usPcFt/NXVUgm4/VOqLL6VxfeFX96u1Si9QkkYTOSdBxqn/qjs3nF
6NMOmlK+hc2tD8vC1FXa+7VJxBUNpIWR2mh8n6oXz0MqKqGkdsea0KPxBNuZo/XAmlBzA/t3lxDS
RV1chsitJEHcCR26anz0Y/qqhW2hzuCPw2udYOL/KbmhRHRaThGK029AsE549P9PNk0glcsJXFB7
3oYZ7lVCmVfURKdj+uX8EMGs9++XZNdeFqk5XOtoKa/UlTTg3t20SwKXy5kPDz22EsNINZnv1KA/
8nDOjc3rSEE6sdCJ0oXIMk7NTEwNPUnSypBlj6rG5+2nN9SsD5qh2xvWonxb1V0VefytSsTFUo8p
BnBHoeI0U8u5kEY+ji/Od/djeSfFgWQP2llW1rMJKf2YZH3imr0t4FuSEvcEOyKrqMpZyK0MPBZ3
C+J8UDfFQrJSOqauWSnEZW1pos5mxJZOxcdvrvQKJ8sK6vClc7UTsyga5OyBso2NtckaIcuRiliZ
CB0VhOZ8jkk/AJkWZ03yHRm79dYSa/+fj5t6f7iCOPjer3oAC089/iW6HftGO4ib9mKdniUyBPO7
ieMIz8+WtV00cOjFNylQUVEh/JG8teM4SE3pYO9fhfXt8/B24pAt7gOUghdQ39qPDUIjvuWZxL40
9zLNjqRYJjdvHCa9p0BaF5LLdd/1oIBxt3Vvoe95mnBITZJk23DFkENSJ3O+Yz0TUVBLa42gDti7
hx9cOGJVwe8M1ys/y9XZdgF6+CIrale/9Ihy136gft25du/NYGcOpg+Uh5XfkL/ugLN3fg0DUehL
hDZU42nS+XFyjoD3SngbTXft4NEWbRw3jgZK7rZ8b1Njl1ceg/5mQDU68oYRcza63VE1GMADyEdm
q8XFP0mY7080ORLzKxupdcjyhvL4qTR0ws144AGqjg3l2zEjTfeAsfaG8iSuZG7/fgFmc+0n/b91
pwbFCV/TP2LJU7qoDTiE1+9MMU+uusbCYl6AxqmOmRtYPbdFbPEutTFabFtdx9VLBD5KHoV9SeHU
XbLY+Bz1qUG8K5lVeTIjNYdGCDNqhzyVw3vsXYP9LJ2zZEWvICGCVxU66uL5DF2LiUB4P5C50d+d
g2u4goeXNWdR1808ReAatA3HJROh7sNSdw66gCG/4lvSpDLH7gvMCz12riEVTy0yzOpTWgFLjLhj
yyaODxLDJKLA/rz0UNfY93cVmio9pVq421aaaw9hz8x5eEaib6FXCOI3m0leFzuuHOVqaupTYcnp
lkC/DvSbuTrG8WYnE57rSPISEHnJmMXmvye/g7aGpOH2CLdAs9Ft+T+zTG+SNVAUX4Yod+yta3y8
tuPXVjhCCd7Dj+LJ+9JeTgSKHqr2XveVXGswZgW85TU3FwASNbuYvgvJ711+FfAkQUulcOplr0p0
Y90uSDk8hAm8l57PuUCflstuCj2eGubulaNjTLueLDcamVYVkmvufLgZkrwaEhAGpm8jUFVWrKsE
rRPwWYw5A83Tg+HPMHDmxpkyRdqguMsU/lCt0tymAPGM3krx0DQhxxuf40iZiSfUT15VDyggK9tS
oEmkD1k47y9i2CVQ6U7IqrcRkyogXxpSjyL+h1J5T8hpi4IhhBTv9D70VXNL925opZEyQLARspTS
lNuMqVOf3DoUVmkKBvuJAxwjArD1H3ffVC+OvNNmGSCnhu41nCHzs75oGATFqyBHbRRKyCduCwOm
RB7v9LkM4M4t+ekYSjWERBrSme5bCjRoKx/IFX42YhdEfQv2mRF/4LMzzl02dFHBrJ/ZN1WtdplY
mJyqLHkWPVFAqPxoWI4BmSi9hu+WhG+MS4FjMy1PolEJOKx9Q65i2g/1MbnEhPIFeCwJkqLKe3+h
0UrOzLrf77EDdBAplYTUJzHHRmvg3N/hbdmlFCnxxLuNV2AhQXNlhiRIg1XBp6lKfKh1vSC8pEBP
VhYitL0yNKgS9sXBgs0+7Lkz0/U34mV+Cq+Yxbrzzm/09xEhu5XVUyEyANwLR2dTd7TTjMHf8nBr
PS9DbHwE/Wv2bFTSTRoyCUfC1BdfEE/pI8nCnDg6az38dziwMvZcAOYcyuht+uQyzeULBRH/gYPJ
riJvt1txyzwjgV1U5hSjYf7H+0nihJYCMktV2QouMcjlTnP4KYcpvBz3Xw9iZdN7MhtH8AwNKkZt
k4wtB88k/Z1JHjdiVjPieBmK9I6vrMec1EYRgAq5hnNKI//YB2YIfOiRFkP6yg7tvRkLB+w5M1Mv
oZBGHk175uWezSQn5uSTQ7U9WiJsfJQpMtheuKaybi/QDmV2DlqZ6XNYdffAFb5tcVAihCyuhJSz
F5vvCE4oi2gvU7msz0Ct83X+h+0qe4Z/6trPRBBfU6YUfr0ziFRXVRLrgoNBDsTzkes5grQ9lP9E
bgdYX5GfDJqN1QpftYKHcJ/HfRJ0P+2KXdTc2FyoiXFNhF2HPrsYc5E1M/XCi0l2vkvZ6HEx9mWU
7vuy7oyT71N3zKX9Pe7eEZQRHVBnM8ZB6+aTz8ts7yeY6mrGMC1rbsDinVpMNi8mcnYPAbAAtzcl
YnuR0xPHFX3vu5Fzqm+z1N1dSLFq+66nYoBmRDrMVNQ4SoaVUnAI9jAJYx+6R1Saq9qmLn5W1HVI
KLdBPFCfMu/g14X+s/yZQKY9SXEZS2VRLihaEm5D4+yEnGVy9aK6pE2L1eLQ3/WXLH2M1OuKjK1Q
cw3EE1zg50hYJzhtryFNQlCz/KtOyokq8NFZNAiUXJMxR1dKplvm91ix93KrJwCcJqCwO+ar7yle
PgR8949Ad7rtSCWyk46M9/PXGqMDbpyJgwNQsTotsPkViE3DbQoVfs8R3WIBlfY6faLUPX29kqZw
85uTQqfXEI+7tf5NXwxnw5jHtAFLTH/ssJwh9Lg4FDOmFE5yYFZzj1UwfcChWsezmuavadjTnyXI
+UJDlHN5dL5lV9qkmA9fp11tp1A1K4XrMsxgScRQ6yKP4djBCTdn8/xHBYZp/GUczXbvBc9d7YDb
e/5xZ2ngPPWiR3RD7KQWFBTUXI8PAjYLNYjYxKN/h//QurGn3lQuPCFYBIIYmFIYqPAm/milRQbK
rTe6XqH8F8fFL0DH+cBlUsVMOIHNa1WGlHgbJPnNv0WfYWXGiBK+MM345mzZ5KLbopTHhG7SJH/x
TbsI3OIYntndZeYeUk6cXLXswQx+yCyEXFNhg21mkUumpuzbf87sm2KNGvvAy4zgOtm3FSIWtqoc
ofTTv8pt2ApU9CWCMPeRpNO6WbPd+5kF9FegOB4rc4zS1kknkD2HiuBkbCO3qs4N67Ai6cIRB6tg
h5jGuwvj+ZEoiF0eSHlaiUyIiNAbEQ4IH9k5BBHkEgLROUMrtnSprJuZPl4PA9jxvHrS1FPAO0xJ
t998giL7bSb40rDJqGyu57vT0ZWz4MLs6SBUTkHvBtuV4uZdcA/RkbOy7yo/ghRDc4HUjTJjIkgo
DO+2lU8RMJUT0cw8B0dtGHnKWawx3/zkJqbXGNdRz9X+/f0a4Iad6HbvBI4yrEO7dAm5Fjzxpto1
PrXIbLwQTzRPxM6DBNR7gJ8K8uO/UPDDnRDx21ykzdfbP/YLwjz+6q8Sr0/V53YlnnlsykbVsJzr
HWeBjjSmhJhlFqxDZu/fD/uXanK4CE2l1DrRCg43L+faPNrBrUI0jYC3lbMVa6X78MJXDDm+bnS9
4EaPMrzhfF72/4yYG/lBKOT+xgzi6+hCN2EMmo8mV4mpMNX7XgHH1oMAAN4kAQ2PyZAvJ95JTr2k
wgUWQj8ANJ2tBnD0YisiQvPbEd3kWbi56RhS6kV1IaErdy84h7nxqrnwKQm+dLb6StPOuWRDBBI0
pdwte5szed59tVFqhZC7L4awcpIto3SVJb7TCqMw5f+Mbr3o5B58e9r8jNYlPpbprZfEbHKSTW9U
GQmCKCUhkMOdM1WnX59zcpgKalJP+qPVUPFuE7OzoydO1I51gS4hBTphZS+bnHN5Jli3DNot9a+b
pO9NsNUr7FIOzaSwuZXWQMmjlObMGnuAW6lhNjET+KwjRhdvfx/kj4VVVItECKV+xVn1PwBkcGTq
0aijY7wHrL4uKzBnAY6hcje6F9+cmb/YaDyN3neMw+6X6ENKSheKMpbCeUAZ9vjYH6/9cjPtfZrA
SJDQP90gwN1kWq+ptCk3LcyJLAOBqK6HHcA5SuJtuXSxJi1OoNvYGVgocq+1fM3uuMxa7B+QHKi8
gWZRBCpyEFDvXfm9pMFeo+IfSlUuzkJBQbxyL/koM1zuAP8fofuThCCyd8m2748grwSAsEZvWqpb
sfX7zygbesKQ1CEdWrBpcQepyYlAdbcFVcCK/TecUU3W/rntY/R0LNNe8zNu0qJll08G28F0edir
OqsIFkiIoqy7UxkEV1g+0pb7+mkIb3SbFbFGIfBlPimoweJQN4Bu0V5LHM5G72+v4momaEUXL7kZ
uTBJtphsLotDiuHnIpzj5cqShKKZIYN9hLG6/PTGB5QbgGgIuVNnen5YiAbQjVpLPwBxKqh9Sqox
VwCF7c18MId1T7rrohSZ9ygKVx1Lol2ZC24+y1C45sl/PEh8SmgHwY2e4rbkdjF2eYjbSoqyquIo
KJP5CY+vS/sLXr65PAPC8PjbuhspLDaqTHIjf7iEw0arqEbcMCYn4NfpYT2KiduGvZ1zC2zrDNGo
t5wqEGAS63z2gQyezrYdlsVbhCsfvmOssiQj/VeCCnmkAryp8V68kQUr+DTru3afhp2XMRUpi2ze
mDZiVTj3ZC95xLQxZjkizHIlFe/sCYK4pFT0y9sUOGOIYe1TbSU8YLehu2ODAuAlWgybyCAWpTnH
JsthKm7Lr/YJHvpHeLpSmACmpu7ej4OZeP3KNjVY9ftpkAKm6KDue5KDlTuzrdwIbV5O/dc/9D8D
cVduKhWMTV+kLWLOGCI3gkrX2+u0X0tRvxK5krzwC2nNxb++zFHmYjpsdUx81VHJRkhcZlQA6B/6
y6o8v5PdRegVdPzgMrYFqcN4n0mRVJmNBI/A+mwaQCnSiXgedyWO+00AVkNpJDxio/zrSCNhZC9t
Kbi51/RtehsssCon4O1aoAfjC6mpT/VUSCfihfvD+guOsg2WCx0S/LrZzPtxDsM8ugKsInDEviH1
DHvOh16GEnsrKMDygGe+jW+8GVxkFwIbbswFiVziA2zAxbPEJtq3pa17R+VxyPROr60OE5XOI/kO
O54LppJrfb6RhUFrEM2gEwjRgG1j8TzWvuDHKpZnG8LvL9pmUY1YmTXx6KRgF7Q9P1nExrICx9Bn
zD1fOKkb8vkKxYdeQjXiRYYvut5zWT3O2K8/N53wo/yXxQ6yL5+6nVVGALQR2Y6sbBbjEJqIl4yQ
9GxqtjCmc9HAVEW+kfPdjp5K+q5+lDvP3t6zL5ldT4N/fZZCnDZv6p4y1l4BZhtN8JmacV6mkm6j
d4m1HfL/PioYyJrq7H0h+TQCBs/oCdyGXFOr/lFL+mM/NmdSD1/uHTusjfBRcUKjtlizDE5FTCvY
Q5PRbbENnu5uZLKbfKyV7UfRlbBXgeg25d1Kqu6WlVGgmlAo4pTj27e6NpqbuA8In1/vGMpofcn1
jPQNg+t82RNY0ObPrfnE2wbT/2LZEqwaDf44yqZoygObDDieQ2aqmlrQ7WqVY5GP9xZrW8368opH
HATUKRAkq6SRLRoIFZAx2yzpDYX+uaQQYRdSOb1W22hRRNfn7Z8ZBtllV2OpzUA0yYqnMxpsU74H
hpcfRIilqffnV3wzE1AvBQn2Fp/10Wi3lsFGLArTAUKIJyv1xQL3NKi9AXxoDDhOCtkJHDsn2SP/
2BkL7hpVgYm5dgvZs1YZ2G65ZPn1kss/9HrNDUuNAFg+TwKIW41XakNVvql2yeiJvga6Wc5WglGg
pWqQNuUeWh29tJIlvOrkx2MiOiO/nBdcF5wop9tBcMRkpipmPDz2AHoZQfvTEcU9Qy2ymdLUWznf
0q3Bzek19q8O/eM4VDNyOVYGLSIUK0Q/kQxFJ8zcjvESZA1rELoGCjVKj6oscW3+eBMBmjZAzEGz
v9+KMHOUcYluhnC4xqUr8kD7pFbiohVllT/kvRFumUf+p24aQQCmljM9hggofuJ/eZPklAQy8df8
oaGsZ6c2WnPdGFlZKlDTezslsP5egRjLzp/x3d+c/jeBR0c3kWoETlpi3/K96vdc1XRGe7Nc7L3w
hpKf9e0v1N1Ut59ESbdpVVrm2OEeNvGdC216HH+6/L/kyDv1PSnOFrKGptNS/m5ZJiHPKObP4rRX
ts4uuYXCMSlGBmBe7Zaq73bxEYW7hXxkgclqkR4kFiTwDyOi3yfdjAvpd/ZZ9u8j4hTf+yBSbNDS
tFLZh9Wa41ZDOD1Y5/HS3wM5P2wkb6XMICdd1h7vpZ4Zs2DymzOWNAYQ0C1zpHaBIRw23RPvGxYh
qy8MihYPZNkMwZJXYS4xSwt2tovztws8LKwi0OR6Esk5qDYB4Gr6/dIP9AGTi/F8YlTBh6Ruxyqn
GTSf/FbCv0XzS6YjwQkHCL4SK/yCUcChkCXvPnye6z4HhSfMJRPdbbXzCzhlzcldzle71iVRvup5
G1XEy9EGSFtDhJV3aRXMt9B/y44JUkuIm17p9j+u8/ZfH957BmsmA/HKZwRDRhj0Q9plf8RCafXV
6uJAdD/9gfRVVRqF4UqSVPzH2/nIy/p4X1dSAPZyhVAs5S4PAxW/i99BaQoDse3XdrxmGwjCxImM
luDsmLRYlSDUAYFgLMiWBkkkbIlbgw7qoOuPYcuwykZ/H3UVXiRIHBHY3aXSUsZjf2aOl37yocpb
zH38yh4XNsR51lnR9B1cnTJWn/+RtL9Yg7BlKb24aEVsNbkcZfi+QJ4AxoEUpwhrEuY+mlCRg96u
DNsRuXk/oc32Ru9J1zSThRtlk/i+xz4BONvul2jf8vDrTjdjMVm5b2kDGTo21LdcI6FzeFusFL7z
Q+7A9N2CRQZEhqQ4wZQNcW6meYivLrp2jQ9epgu5Vwe9jYtyMRf59JJf+UFgYMWaGrgA8L3nQIT4
jcA11G4fNADGeTmuQZv45vsYQ4XgwmIuWfWde/sAaswuELbwFNNcIuyabhNMquBaxyHvcK5UwkbY
7oZJyhfaCxFdsP746pZC8WLhJgwSMLZQCRJxaTuhFOUYXl41qpqIIrwhvnb44fWJFR5usE72Z1pp
vENVpNIFhxzVQ+R7A8Yq18fRq5M4v5RduOWPCwdZbhNYQQ35bbhp9Gv6HSfnicBDTXmpIpIDbeVL
CCr3hP7OUIvvpsqgDi3DE+Ud40ldf7Yk0RE5732AJJDTafa6GivS8UZTNFSW8XAdPbyoSP5CDyw7
oxMZ9p98kd6fxJflgSRvKoPTqkPLzN2r3A1+/8y0Bd+QAUrRLXh2j9PUSzLxfx6stiryNGVf7Txn
ibv5iclXTDsZID86awIn/aqV9UrIbV4oOOzBdkKGg2cP1RvrGmkqOyICtYIyyi0G3h3e1oFDxP5Y
/Aj3i7vO12YT6aVGtJUM8931IkI2RStKM7HUkiUKb91c2HIzna6nN0G1GCl/F0uHZNm7o+WtYK86
vr/ukIZOCdbQlhG1ISyawH7WDEC4PJMbEJYlci89ntvURAQYUTsFpauCm29rNbGLgEBCql/48n4Q
YPZOL2GiJvf0RO7VULr6tQxPmCNZCthQ7ze/aghh1xzEeu4ypZ1rLIO3zlNb2kSG33rnZtX7LD3O
HMlMGU7soVhU73ymBIc8AdzgxsxZ6Mi6hgOApIDfRTymwLLSDqqJqc8TLLbyZeIBJMHVys6I5Pal
txFcpQ0aO4ZMxi7/JQQQu+n5sDFbbt60eCcKcYA1dfboC7qf/KhddrlTxlWINtgdiaEa0HNFymGc
cicdmislspi30T5S/8ATf1Y3tszCBMkc8K3hNx/qe51fZYHW4RjCABqFP215b8rTgUy5L62iHQ1B
ZyWQSJkzKNzwYezW/eTenOswHkQhvv3jl7jGgUHUDhJ8Rbu5XofPmtDxHZbQPrfe1PcK1w8rOg2d
4bDe4TwDAnIWeq6kNNQE6lED5QfaDkynkug3C2fTNbG5xMw/9JEQs7IdLSMmqGAt0RX+7ghEmxrM
pyDJT0wbnsgqsz5V9IlHNhLzfLUv3w48BYwjoo4lE41FjVrcWedL+xQDHJa3zUgE56BHYdnpUFAs
Hzc0r1u1aLae4LrPmlIGxm5vZjbaCSjg5QBT6joNdtRb7N1+ctSuJ72OrTXy9Y9l37bhRQjuqDWs
MShgfKecaLlnG0uvvJIXlGITkn22JF9hbL31gH9N5DVqLP4i02HQVZcjEC6BmA6yRyPM9n4/6tLk
56fFpLmgvPta1w3ayliKItc1CleTp7mhnziMC4FITEjQ/cJAKjNVnvHerFZrT2TkV/eOo+KKunJ5
7l3j48XtHWb7xq/HWHT22zuZB8Y1MglO0vIofxfq1eJ5qMSkW3PE+oEC2Fmy/cH4u2ABVHbDwonK
lsK53SBw0uuS6UuTePzrHeBr9ArDYg/BLk37qP9qmsOwKPTCtPblz9Jt2uELSFa5hDWlQ80PpzhB
x/kmxEJ5RQsVXI1JGNZ5nrJsDKMkhfmpA0EZ+5Xib3/ehBGgobwRYM0xuhslze4IZL6mIa5U7/wX
NewPrWrRk4Zo2+Bz40C4WzBIouikM/2rTqOD41uNjjLDvfP2e+0chIL1BotggP9TkkKKNDgUm3OA
YjKh/WUBSYk0u0Wz783iA480lshJ4b+aJrFMzAQpckJCTGrVbQ5QH5ogpe+QJE0h1IqPeRb1SN90
BywP2lJsIlUDtdx0VDtnNfCs+uZ/EUMwXjCgoKcA5xaaF6MSk9NHb9FBqbW5EaGnQjHWI+M+9rWz
dcTfuheNc1ZP5ew9W9gUQQWzb6eDSgD2cpNFsO3fIdkTS79e7yfiZIidzHYmy/UWLwhN+3N4o8il
17MHR4BhQczVnYlJiMz96G/z7Yz7oPP11nNTeW4vEVdqi3cTXb37fRFq8UF1qCGzBSyZQktkBQ5O
Hp6fg+1iV5jxI/jcNshHBsfK0NpLx15e0DjatnmEdiuPo1mElTwx+/obkLVrWilLdipTNMhVwa7h
uzD4SggNa29B5SLsXYCOc53fmimI/+k2pHGio4j8zt8AF1/rTacZ0OitmuE+lmqXCB+TF9fRVnQu
KQUJQ3r7312BcxbSNk6co33qYrhYNY3jXEbe3dHw4nsUj2zheQkWvEOzFqRsLk4TBNPjoS0+vugp
oj3eQRpiejU+pxqzronBd8thP+PfWrLEeD4mxOxoALBWW4QsK6OXFLLNH9vgbujOQuvXCIUkFQr6
3W2s8hXDYUx+XA81JFmyWrwdQmE236i0Vr2RnE/M9iqrYqtfVnEStmMftHgdOLfDGHmtJ5L872Zs
GpMNMBTFwgGuOhs1zZi25ObEq1Lw4SNQGVzCwC1qWynbTOTdJY7DMQpo+/4BiPlxHLRwvkJ1kI+z
+/9IBW+UaF2lMYH3lOTJUvmnLib33Z7JsuKdyaA5dAPFlKxW6sUtyjcIP2ayX6aka3z0Nyr3PU4c
aFbgqZZ9JDrLx5O0NiG1a3P24pVjIsEQuhDonuKYRX2izMwRjpdpdky1s+nZl+9f3YHPVeDHVLeZ
LM1laAgi2C5eGa8FauH9ETyPI4zxz6aci+3ky2q/hTBniHNnG0HBPDQSX6u66Ke/wHzoJV0DTRoG
7hybcf742LFRCq8DRn2nlbXUPlcIfDYQOxulf72/JZnqaesspxmZrw+QC1FxbBxXOm2OG6HjOXeI
KNLQVJ9Ap03TONteP8pPJ5NUC4XqnD+9FBfyAGoXMeKWqqCirGxCBQ+zSouglS0OWrSXTW2hKYBF
RtUZJxvbAkEQB8gHAe1KRkph99Xbvna0DmYRNPj8Vnd2aY1gjOvQMWoojg5IqLE2HXHWeGYs/bXk
aqgaBgvtSpbMRVS29bJ48tTusGB8nStPeO5EBO34UeALiJJ3WuqJOMI2WfjmYAbgOZDoD7fIplF6
ZeJfApZwO0Ix1BfQiEmwLAXHFVdslG723PaUdNXJXRhKkqjkclEi/lmbrUoZqnSaVFY/Zs2OMF+Z
rFzIByw1T72TvfoIsdRoE0VU/ZJClfjs1ceP4Iwjo2R/i1ZPd7ZYt9sOa/YwyATdWWTgVVTaCeYj
SIo3kProG9zbXyKNfTyphOsSeB6FVhjst9kbA+fE5Tz28/Dm+vFr9nSqh4gXKEYlYWMiaF1vR1yh
rvwBrpMfITQ2Y9ouBIbF98mYE2I9xP03NbEDiOuLjooAnmHrHG0CMtkoXeVQw6dTEndP2e5z1EV7
bXIKuY/N6wlzWXG4+cE7fGEQFuQU73kTsJaa2V9+z/BnDOOJ9HfYeMtDiEdRMuTo6cgkKHSG+tC9
AZ3AzjgETo6OkUFMT8pv4lLLp/rzQkJIwmz3pMLkvNLKZMszZ6bDQmF04gvIn9JinyRGCtOG4iT5
Jw35pjuV1rMKKqgq/wFX7P3c4uQ38qwPZf9+kB/U9XUXzhC2fauw2ltXrZm/dYrU+2TN4+TOpvWL
ChYQXN1AQyu+INtI/V3VhixWkURwXNdHk9xsz9Jl7OyepzaKlSKJyHSmloZZgN6VT1u/KcqfycWL
OiVTYsK52tQ+ZqrknOHT1MivwKs+GzGKTx1A1e/9mihVibwqvb7QJEuPwU1k4PPfVwVKEFqae9GU
eo3ztepHGaT0MQ8TpShsMet83kdIE+PqGWgTD/j7VXs//3gnvz3/MlJKKS/Lhnkm5Z1Tngg29M7C
tqBkGyexHbxC43yDVH8S2rPPPKm9KuuPKrphyK+4dkC6Ds9jcNBiPZo40+6FriMvFe5S3qZmZch3
lHZoaJapcPLVCkR1NG63ejULHeRWOJ6GmNUBnFvlGYdg4rsw+wQlI5J5lX2XjEjVFik3sSHdgRiy
PY6OJfvKZVn9IMOqoD0QIwTcf7jHXTpbagOu4GiWKsIUxIcFD1EP7Sk1nMplLtpcDsPMf43pa92t
4KW3lzpkX0VaW+K1dX+gJC8GKhwF4D4WfRPHEJ+Z9+tpq0qcrXAu2oFzPNmZ0tonL3ogDMiuHCRd
4jppDnWkhIgOuJ/TGbBR+YW924FjPdcMK3y3NJDQDWeGVE04wSixaMiyYTiE5I7O2lZBwsTnvWTp
owzc3ynSxxdpg69oOg1Xs0t9LmyzRq5D4/ISw/fJr1G58Z69pp8rJfSbkkoRU8opkmwtIAg7c3LW
ptmIavo73RzY9qSKtXsUQPvceoU4kFQNgsVw/pnhJPDl7AkpsJDBUoblozgtTCXH+Gl/WkHPagmN
czEZWM8JziZLBTGQK0E5Z3ycSb5MCorbjRwcP0pqEz8MMLXxxO/5EOMbpfD47w+cTKQkcrX8svCU
gFthPXsikC7F+iTr4tNXWorPVw3bwGfMxIxv/4iz5j15W2XqUFZ82cy15bJ+MscN8l+35xljF5Mt
b2LMUd/Sgw+hQloY4jMeFqFg31k3Fo+5qp6udCSEN+rGQXgFK3EIUy44rxrE2+2xIwszyW+25BMw
Imwt5xPOsY2CvQO8IWnIcKKPZGRnOJoq29jy2266DSWhMvnSITElEBuqcf3vyzrD/8DZ2oil8xhx
M6NyTvKz3IDnmGPwOEw2W/P+ufKnlvf6BpjBY4Ljs800TJyfJJyYzr+XtZIOwhiHFyvjaahyG6zs
0NL/j8HYVx5WYAs1RjtwkHl/ZEzMoaxcFrNNsIoOk2u0saZHnHdGYAaeVfpO9TJ+FbX4E+gmep89
5JONxzqay+O2zmYXyn76GrYKofQZ89eq+6gOQJOrm28EUiwqFUprHum1pFDTOm8UpkysZgUCk+QZ
mVOVsUPSM54cbYu/ofaBVEKpXIqCyisMU4lWpzNnOEQo8Ez0qpbace7e1abdrjeaQCF6SOzz48Cg
KDyP5IRitCborJfzZ1J3rP793vwa+ROkRNi9ZVYPGPldlZbjKFLe9huGxB20oijLY5V8J7Dy/8CI
Scti9tlHJtDLF8M4jibbAywCnjFYFEp//RqCcYwk47RXdKo1oxLmPeROJRAC1s5G3kukX4wFzXop
blzhtyJVMYrAe7kRdcYm1+vbLTnXkUa3PIXEr0OtetmlaBPZlk+Jqv92Dh48uJniYwdqZT2LUBLa
xNWp+oFrdIWVpjckM6+Q0h6QJY3gn1vU9GpJkvF9AVDmY4upxiCVOstwN4q797e9/+l2Q95rHT7P
ENSMO4x8WFVKkdlJJmv2izd9PIOnPDSivsWCCuFt6PNmqNzq0lF80xPD6VRHgXXUHSH/75uMtIVM
Y0g2cPLznB2DzmXi8xed+uSdEa+h3Uz9ioIS1BaVUsXR3TOf+seT4a9QZdzIX7uVmn6NP7UKkaOU
uHuUKZtn/wuM7K2YsNRbeeMkjU7EQ/mnoSaVL/g+RzeD5HCEPyu04+ea0jV/dEne+EAboDRo4h7l
p3w8e+gC1CJ6oW6+P9bEDlYSKmagik0kJXZZsFIsSwm2bF0QCbkdfbd9Qw2Vyvop4FcKttBDcaMX
Wk6/v+uWz+h2iiieNy/Ja6UwSmpPSKK/ICB2ZIYgoEKyty966Q0rYMi+aFAvJZpSDJL0CKq7TpVs
PUxB/nIT01P9zIXBGa+4ZEhPnfhbwRJZgRFbc1BllEU5bk7Q/ycV43VlpNQo/OA90hvhYbvVyCBL
a8dFOAii008ZFaStIXev8DEFUGpGSpweBczkxdgxSD8cecQ72AhbVHRTVwZRgt7DOEvqgaflSjEn
niem23hi8dOLKif5JhpBzRXaSMqLdInulCGuz5kSjZp5ADG7wKM3uYwF3yCHUnmmCAhxwIzpdDcH
QVmR3042MyU6M2ptoSviIaUXoZEcuqfhzrc9WerHfJ4em/eW4B7dHixR6en3UBPm+9jBfOPj1BZc
3uX5dEi8HEkrxaWtssSkI/4JIkafox5+ubMqLj7JdalT0SC80/k7OxZXHEgTrfvUdfGDlUh25rnv
elQVdAAD5NXDrXyRO0/7DPITFnu0sRXRcwCKZo17MqZ9MPDbDNeVNibMVcsTKGHZOia0TFMMpGaM
hvJ/vovxPbhFMXZCiI8kr2JDkj3XiLQU/q82X1ts4u4xsjwtKWrpCgF/iD5cYqnB5lkwMGhx3J7j
XYBAG2n/ayF+jBkok4+0xBCdtyxWKOK3IrhudXPwfASA77PiK+MyyTsoNr9Oet0+8vAU8/ubOf8V
Ft/eO59j2D5cxn2DYXd/R2tc0pEQ3Baxz6Xta45p3Qkjc6Ul5JQLd9pWq/rKqRGd3P7moxqxT/In
fYsTxtMUYL7BmGMtm6A4IJ/dzm5ldkubV+WEi8atc5TJ8YFjbNG7dOCqPUb5wtSZzNguU6ura5rz
3yg7r7o+PfYF2vNlV5SLyr2qapTOVSFGxAHOI4oVPZijvwWZrPGm9veuEA+DKtmzNl0MCc6SX4mk
+zNaafmVo0E6R1zXAst2SJncZVTTjxZK/Gu/uNSWVb3GZaSyxEMzrPwAIkvpjMMrqY8Ib4jBt48s
OCHD6YoX3wjQTZG64UHp/iJaAfxbwzX5GjPFSvmwXdtAPwDo9d90YEDzrcXaf7dpCVRfQspDRMKt
oa0kU/PAnWqVkdyX+bq3wP0KB5RUrjM4rCiLxuxWwh7mBg1vyiVO045oNOmA7AQq2tmkujf7Ww51
wfPhA8LBBh3MzAa25qo4YZMUzG1W+5Ej66WDd5z/o6VrGVgEajnCrnaprxv1RbWH8iBpVWqlVdL5
Wvmj1JY0vrJe2MAAwMZ9GaFxYiuoJA3AOotaZCKyr3yeszlyxVERcO/cTroYDpuyFRMTlaF3JfEE
o/UO+FbvFQN+SMaKU5/9RTapIg6q2nd2E1V9ImmK4JI11GogkIoFAPSZYHTrUleI8IpqudQgTq3d
uqyxwV1QflqUvFGdAhTzjAVPIGJua+2RK+JM6rgi1kx7jxr+UOlAs903qAe3xWgton2FsG7OXMh9
QAAQCz83tR9MMl9izsQlEY8tYeoqe8RMktdCBNCfzZQ4N3LjmLpyaFZtOpD+XGVyMpaqdG4VF2jA
0gejFU/hrRUwXDZob1ObD10cZ5OpNnqK4tqMMMKKNUh3COsITBkQLpX3c8Bh/ZmuMl2w7bfiAr43
IWkdzD08fM7IW2cUmWVqWSdhNBY33tgbVKsJRuKluTS+2+L1hqSCpFhs+NiNs8bJjG/iy+LVLke6
SiMwixI9LDbgJbvyFW2eCo5zJbNlWEvXouqPxWQH2t2hT3crdEdu+Vts6C2uUbpe21z0zYwKExdL
pQxGE/ON6FHKmzktie63BWiGR68z73wl/tq71CxwcdFx72O06aV4anO+8e6wUtaYesaFzB9lqDE/
eTowapqOZZLmaMe8iGn+uextamW7MlIxoNHiIqKnjLUqqGJi2uJyTVRemzJ+Y8jbUbu13DqeI75K
g6ku3GxYwi/SmJK859QiBATJ040RFlZtoTzqeRuJ7gKdS8del8iYI3WFIUDnYPcETpIPaSV7CqKT
QVCV8ivH99S5d5zmi6XiuYLU5DQW4LyrNotAyHAKWrnYLgvpUZtTfrgRN1pnm0iJ7aaLgnRr1nNc
k+UABDOtMWqiphAXLJgxsEDSw6wTndzWPYtHEcCEHK4yICm3cJC6V8p1cUbCSBcOsHJ7eBua9X64
fWa0gITmKPGHmZ05cnG+XK8ACkHXNg/MXesAVmjZ2zyUhXk4ab+ooXeGKiyCeCETFzACXWRjjg0V
DMXqJx2haVE1Mffw53UZd+lNfWqpE7RQQLa3bdyncvG/ihkDXLYjPkMsGihQH6gQPXwkjsbliohe
QPi3jy+/r0IRIn3DW507O3XAz/U08oPHUSgWpcG8cZ3Y7oGB8Px42g7H5DulotezK0R8k81OX81o
02le0AR7lUqq3qXcqJxQxdsJ86F7IA94XHd+EDJwPLonGrjx15VAkAN6+Qs2IoJ+1PhMwJltPu9I
pe4Cujv+O6UQE8fcICjvtLzEIJZ274ZB4eplr521AkuRY+SVwN69pX8JufNlahfwlQ7L1MvwkMK/
JI+LPflIZepbijp2HwVr+khzyyb8kRWrnpt4GSzgMcjmnxUwo6of2ssZn++jvW5uHmxl1PyWnO3r
xBuljmVwWzhEN/sWLtulZgSRAFhpU8qW9m1OAs2A5biGYMPXCL45icZea+2p+ndeUyZ7QAGVAJDI
F4PtewD15J9ogNSiQBcTsf3CU05sRdz1FjNcKdbMqn6irXiRnmg+MRGXKeAOr0lt/x6VxU/lLOMX
XXGd495H9vNHf0K0H2QjWI7TcPHZDd0E5+i/6c7MzZEWweQFCC7jhZwz4hUf8LezkCpHeSvbiFaI
AFWExRvrLCUwJYEFgrBSqQrVIbRmzIuwz64BLjmikHFkf97so3v2NbVHgOSUlC8g//J+56P8UD7F
kjz3Ym5eEIsqkpEZiH5xcfdk2so3AUEOc8AEkbPO+5IPOv+o0R4H7J/glq0BX9fS5GFc7bG7nIEm
++TVivy2UakuyF+zV5xaPcrqLzJpA05QhLDOxruCBCRAAMIXXrRk33gCb+xVhGPwWzmtE6bZdGsi
ipYplZ9GHiNY6dOUIAcCCL+5CXH+/AWjDZJfrToUvywEGpHBX/5ADP0kGDn1tmIA+z/OPWieQf31
CPlfyLn9wDw6S6+V/OIbPsBJCaMNF7X9TOnXjuXVIUjm2Ph7bBesHvxYsAX9Yl433maRqfpdJI7L
aNouT0FIISEgbr9NIPJb9LMWUGYIWniP4pdjLboou2I8j+zlJLNS/QfKQBAzdrAXm54G5zmqDY2z
u62JbOjSq9nhRjXQiI0ZpRoj0bgZxGKquFI3pF6Vy/bLk2qSOIol8a9BVUHj74wTonjnjBiOb92L
GsxjBDW/FuhLs9Ncv4rXTZ62dhOl/J/ZegM1UW+kW9I0ARtoG5K9h5IRR1+4uY3603uBDICRNIfW
Vl4xAS7xgJykN2MJECsSvdheECNZrrNMLhYeyi+BxQUB655745o+iBEvnU1h916vmuPYZ+AQyYjU
y1qUNgu0AMFewacMuGKAEsfbFKQ6WtdlC5YQOXkVBQ72EeCbG8OO1+eZXbhbMP9y4leN3XezGtX8
KcTLOXaQJK3C08TjbDmJUVr2sYbb2iXb4tsePIG0iGcbGkPBRufEiN/ZZ7z1Lgp6rR20wv3G3Awn
E3bJ6MbTo0nNI2Sno8hryt466VmvZcUEOQpK2Gid0XKIFyii1TYcrCUE1RS4b8bHwaI9AzLExqje
tMdotyPFm1c0LYmlIf0WuSAeQ5qaQBwMMCNhmc/pjzV+Nv1pN3SsQbglRCwqdhfwyHvsGv3FxdLB
w/rD+ORIK20wI6cE8gAwKrGcJdJ948SQinlg0HrkhebQWUWdX92siaMkC8Zki2fJYuNefp7QduVM
sU9t/nzbhZtZYqzxbBNARLtNukSWQr/a8I6FtmsMtzqzeg9zk6wPllbGQjDHNprE7O3ozp1gUZ5q
CCE+q+k1bVZ264LpflhTKPlacSJ+Kl2I5QeVI5D8gR7bHz6gVLk/IIHOSFjMEpeOcu+BkBG5s+Ji
R+QudwD3bUD9aqMBLPmVifZh3EWg0SPPE97ESl6+4kvuVK6zFz1Uc8Z9/DT0ssYZg3B3LQdfNgBl
UpddEvhCsKCTShZ4uTZt80LzPRaYSj/LBw09UyRYnkXaEgQW5QZe8fawQy9vznykoG95E5hIEQxI
cdvLo4llOhF4BS+AgmUS4O/wPImZLj0/hxBjB1uY6sexnrHckcQUAvNz8HP+NjKbESLTBpUgLTmb
gQREJIK8xzLXkrdsxKQBMH4kXCFKlh5QGNE3omas9g7J2ny7m6h3yQqIpePmo/djUR/x/ONrcaSv
mFqJnOjizPV84uvV6ewSqXVyebX2cH19nIgQkeBJVPmrisP+0Uj7dXNrCsm7AuzAlU+Vz/Wpb0sP
ah1CGprzxbzIjWnbxAumpfEtM+xSQRpTvj62EpSpN9vHcESmxjhndju1r+qLztvxOInC1+sEUuwY
/NNhayUNBM30fDYR6LQ4Otfj/qfsfUekFw0WxtfAY4aQOp/ur37S5XjzzIjBQxHyfBuSNo9IeybG
4Ai0/An/bV7hjCqS7oBUOz68wi/RRcrJQJtXOqpWGy0reAXWjtN3iVG7hnEJ4ZqykuMpGzuTgbj7
9cpEFDmsxh55LKp8d1A1RYyZCLvIBREsrfBIMf6LwTylsTmm0WVTOJb8ieNaLRKP+kJvRj50Ou3M
LdPGBo4LC+GXMX0VuuaW/gDFOZ6PNFUa5W6ApW4yXeJXDNmOjQBtNC7u28Ebw823u4Tfz4fLyVFe
l7oz8AvUwU5x5LgRhI1jJDxDdt3REGTYYOXkUUL664gDG6d4a13oi8l6C1CRYYRMpfZpRuvJuoKY
MvXeBaN60bYPQn87xXu6ggOVgsmJVE1s3fxhUsTFIN887uzrBIOjRIBaVqQLZBQvYG12w3Lg3mUs
I8wfnhXEJ6cUaR9iP6P1zfhSfVZZYzLY8U3zBYp/k+78OMTVe3DUD27pvF3nusNhnVI3Bfb1UMBU
gRvd8EmQKiJs8cHysruOZ0zDhBRuVAki6gUR5UT8x9bNt3K4AfnIA7imnXauAxruSUaNCOiSV2F0
7qfPRrotQJMQ3yESPqf1/xc17KTdjPihyfVFtlnlsqYVgKmJnzTmNzxkcdgbagrdKG1EHFrkE7qo
EDUlyn1a1sOrei/FQemLext4eOa9Xo8FZPTD7OwueQa2rDjksja6vSiB33vy7rzFPxHOUTl9Lt9q
5kp/JKPMOatKMXOHSc8l91nA6CQdFYYeVlVEj1IkXQMfvPbzDTlEMWw5eqntbGtCYNT3OctgUfch
QQhFR4khrnYUeDWUJAvEp/0eNGvAi4nV6AcykmwOsrVIbVyJB6kHyD4C6Wq+pyixmwKDb15JELYC
WCl96NERBATX9Y2sK4hge4+VQUmj9oB64Sw48FKIUup/FpGCoXpQtnVEmKiV4HFXOb2Xvx0lrThp
IyZusKvPZwG60CB+RobD3I4EJWxaOkrnmUsc1asoGa5Yl5S6NI1pjahtEwErrswmi+/7O0QKFBwu
UATQf9RzHQBaxdIw3pfEKD4KveFBLfdSES+5CTr+OA05TxNBBaRRXi7M3kpcVbzUhwzOWYzLbHRB
kWbkNndzeKqWHZZBmM4nLZjx1IgeaXmvk2eZ2FedipZ2krY05K0xZKsrtO6hTdGykjOg57pBgzag
MWGqSIqUUY4MFB98tSd/h3tNnRyUeaX5KXmPRWEsaxDqsQL8Yv2PENh/obAX8vhswuKy1A8tEPgC
TzeHrG+DeFQ3tPyg47suzuYVB0ybH4uVD1+UJMS5rLUvWtd22Qz7EJiCENps0+LjgA2O+EApreOS
nLFeWJZLXQu06Nljs62jz/Mu3TKEeRXesnmDO82HnfDN2YPbqiytOt6rErByzHkjIgwUZnbPPN0s
3I0MwwCvxbn4/VC+gJEqSh+vxwq0noaYBw8DWBjztwMNNsyppH85854nTnEqEL/fdjbUyA581pZw
P8VaX7ShlgUCegzndZ66DcgUiAJlMtq24X83glr2M8TequpslsGmfK3AqETfyNaSO/LVRidfJepS
nCpLkUasFhjP/UXZyBM3bU9nIqLOIm0Sga7ZE3X9R4i8AJ+UNZ/Nw7YfTDVEbvHhI7x1VoBjqV/H
w9NoUkSYyLmVcsS58joklSrNXxuXoRN8gq6i7OXn2hzu6FiyYKf2jILDSz3kFqb13G7qyqy0YhWd
PbYx0lL4qCJYB0rWddDaR8hsTrhe24KI8YwafkkBnlFz3zqaLIjgZYI717Pb0p6aPREt92SkGrbc
tmMc67ormGNM23eL5BCO9fvrsDaSKXiggyrXZW8V77Lg4FA7kEaXVpS1DkSA8hQw6Xg0WwRiFV3J
7JkfO/40h+WwStRf79Rh2HAq4N7CcznBqYoZ5EFDKLDx80QfJKYgO56uz0rr4ADtSGHW9xZgAsI4
veIHCBysvOVE8OsljBSaLVh+1yFsy78UdKq7EM2GX4fUXziBlKIVnSulwE4E3BFqL0GGlCCpEzlk
4LdFOERnktoT8pR7+HTR5FZqZpPWWB+o2ky1hv5B+hqW6zl1J6D+VwK9xJ7Y+589AGFHCpdDzvUS
z07aQzldDzf6raNwn6HlfVqBauZzFcE6LQ79WNyoM4B6K3MpxOL53Y8uj1Lxc1l4K8I+ZwyuWkLt
DrfAoDAMtLu2e9kEmGcR3ilxNbaEM70cwJ+E06wz3gdGpaMMqL1Yn1/FSBD1516b4LiWzIWa0Xwf
ErPjd02N96NhxD00VbpLYqTE5o4eklvXEGnivqG7hbk9ibVj8t9VddtuMeKUJwY3T84jI9K01ze+
4oVh+LZIYm44oT4wZ2FpUNrDTsGpA1jjTcvkUiMhspOMLmt8J4pU+H91kPeKGcSlxleGCaForFTm
RI7/hEnOyt2LSy0hxBZ1GFQXHLUr/oC4Ag6GUztlAq1V6EOR3J7a+JaCrjPBUmrFSGVaBqXXfF5t
N2Wl/CSpl2PqhmnrIUyukFiYZt/ymusJ7tGXZEBl4preYkbEkkELdVWyVoBn9xTH8nxmuHpWjDlf
jvhn2fPmDczTypgvZrFMdrER4WD7GRsFbsBMoyb2tKzxGiv+gw+ENys/e0TpmxcuY0xKsyAom3FZ
Ntp121AYaLMQZX/uRwQEijtPJOvLD+8GFr96wHi/lBlU3/KHhSIRoUcg7SQ1EOAJhskpOkd0Hns/
LL2R6xyE0UDdYMDS2UPfHscK6hr4JTPwG87HwYvZpS/tFA/VUuAvHBBXbvISw4MiEnF3PPZl6fwY
GbdPZB2esMcAJM6kuyYsE/17jkqNDnDH74aj1lxuiuk8xwP12gqnRnSy9tg07NVFkW/v4vPiHJGI
/RKNWyhi8DCLpa8NqFJ6TPQotAMP/3BdmxKs8WXB+XtV8lL794y3f/BM6h9MubBGEyEH0K003Fdq
D4McckOxwKtAcQdPr2zGUBx7xx5SdfGKKfSuicicmmZFxMAE00a1/dDiVAtu9gbsthB/ZtNeq67l
CxSt9BI5cMIKoMjk7WV+vuno8SeTJ4lY0lIpn5vOLDrYdArMonOGJfm0Bq50nmo8k6pYfVq1A8Zz
e/ohWKoTyuXTsCY0fKlLeYnIae9ch/jhcqAs3OhpGw8PvcpEESdqTSh2xpU8PGT2BeJjX3vEJs4+
GkOfqrJxoVjbzLbAUc9pBw+KIKbk8o3C/KVlcS4FVwPph+MHwm9QvxHi48NppO4jUJkjmvdrgULg
RAeCjQ/97nwF84LXV6MLiT90gNv4oF6f/C+42YKdI0wAIoK6kmKAn0veJN4IucQtLvOjScCppAG7
mcJdGLmT4M2c11Qlt6uGvtm2mn8y/14G5HS7OavJtAxLv7X7/4NqLousBu6H0mxlloBof8awYX88
8EqYPU8i+YcQQk02kzeUooJlAPjfp/Pub33m9h2vZpp7sZ55cu/6gGPtcnXoX2SOo1N+2WmwhR0U
gdGtgLBCyz7EYqo/dLlSQs1r4nlZk8JB8NvoYoO0BD6vXVy4fGkDjP8rYnMJgMtPoXtN52jy2nyV
O9CFGM6WcOjGPjMtQ4L14lTUXsw8RrB3wfHuCZ6VZFUN0rlL71c6nqVMSYuly107mQQOSzy29Z2r
7y0zypc+Gv9r/29AwxmSgrWr5DQepkmDDxEVNXS7v/QENDQEFRMx7cAohNQ9OItSkl6QBZqG4ExQ
exOIuA5/5wrOHZh2tHEXsdC6nPUP8yRuEnoEmgkIQvA8Dql5RmxrR99a5coZfSNY6uHPeYTBoWB+
UDBhqVbCgAFhtSgAN4CqMAKXgUbRcObmdheWcrNH/ih3mRZoPQZK/aPe2x1BbzLqF+VG1LkS7JVc
5ioA+5HjcE08HaBpyzkJen7qC99NcXSjDdbX0VDtyqtyb8I25qx406ju9NcUpIr1rk7JoGpgMNTg
LoZufct9RO0QGC4i+PfGcoqQ+phBeDQSIfQCwf5pb1buVdpvoMOgpZ2+Q6WrKjJSuIW78XERinJO
x448pNALCFVt514xRbvNFFPr/Q+RY6ZXaeZ37AfEDNAAClg2knL/pVpdhdO/C6O2vE2dK0QGgmMr
vRT+4Kw+wkxtEEZKGfctAlFQ4zrD93TCO36lhOH7zrd4RK5rbfTUkPoOzgcUC1eBbS2zUSkAZ5Ge
21dh3xcab+3WWYM1ZDBIth/s401Tk0bgGk/Itax/WTUZY1OD3pKqG4XfiXUrX15fysZiTPOtBoQi
nWfPocTKVG44sijplekQRiOxEDd+CfwxY6nw+1K7ihWCg0YH2ZZ0SWbE/mLx1hboTD2jZpRfCkFd
pFefzEsTzVNwkE9463S5ax05i85h2BcWEv9zMrPU63EvwhzDkGLK8iXiwHrc7FZmpo+zHB4TmWnT
GLIM89TvELaTIjwzbrOUkdFBRObVVZCU1yADD+KbbpUV/spcktt3+eDXDLRG4dwV/YIu//9uWQZZ
kQJ1hWOtpjI/6v3iEclNky0QN2n9su3oOtEagevDcZGt2ZbeIMHXnbK+jzkIanlC+TynVaMHlHV+
cjW+KlImC0pxBpfhYRvRdputoA8hOFAYvHN4MUqiQ/7cdMwjGbzdRR5i7OSKoRTVsc1oX6fXDDAS
4KM4/CDJfIOcRcsLftM6U4FOqbioyCZ7oHqc00IZR52WxaumD/9CsWX3W3eyCbWpmf0xrLs9DMSv
2PSJj3ykNzqTWQl70bMmAt125p+qV+0HVP5odaRrjEgB7U8M5AdWUrzuVMChRA1HguVE22R1Ebwd
2DCF3r60xivGBJok7kVNDzPqBaq0Ld7W9wVbusW3A+q9PihnWlmHS/3YsAPoWD17+F5LbTSnwPKl
A23Kf6XHKAU6ITPzxcTlG1mSZvm2vNq7hQlqbEAH3m5Y1I0Qh3pwTR+dDnvan0UaiRZJ07SrYa/a
TkkUTSaRYsguVR03lhF2NQnQogdSoAOgF+rfPZAprjSBqvaKbWgUDyMjn+i4mhMdK7HUZedjcVy7
uSYzGAtYkq4U75bPIt5dR/znSILoA9keg8tt7blrkRSQQVvq44Sdz5N4/X2uKD82CZC/crMvWIWG
1orDiLdtj7pE8+ZfzouGhWFQfxx6HHcO6zCfd0XIKOlkpdr1pBGAX03kRUGxiHW7fpTPdJB0hjFb
+2k9m6apW0R/dbXyFXWrcc5zSjcnVy6XTGSMCFSZpb+Htg/XIIAmglj4FSLQr65q+KlH+j9tAw6X
bLkwCKi3UQ/3rOlIgIWKozGntRku2OVJYZ1AgR243WBRurEny6hxhWCdm8dFMx17pUIE1iEv5/8N
6hsDLQP9na1e1AN8Xy/55kx7JdmKExaw33uHEuiimHv+X96F/rPTM9qRNlVmwVOgLWUcuCZg0+64
H2cLCIUKHWV6DvzPDzNpOXMZy9ibhOuUIyKc3FcqZp+LNhPrhN6XOg2jlHMAMHtpLtFOZSOu5val
mYg8Fc5i72mSKA1lTB7puELqesQM/p33cZLDgzOUsc8fqviPuv0XcDJN1EXLYsSGR8HGSTug2ezw
fPL/waQP6ueMe8Dd2x/GrER+cyeTwmjry7hw0THU6YLqV7Vk9ZQHxedJXbrx/CjYV15pSOG9GSsJ
88+0ok/7U+dVfGywKGZBpgJROBUVgLkISMBfNXmm8bOyxeDTckoZ+niWMhF0NKD+2WD4pYdSUsD2
hMi1qlpGW8K/l2YsEzAH9E8IKxRkoF/w5ZpmZTeUCSvHe/b/6KFNBS8tUV1nG2wp0UBJzhqlgpXL
R7Tdoffznz7gvfT93HVCatb5K4tecf8j12zq5eAQvUDwoDjUqB/PMii1nC8s8RT0sGP13LMa0EJ/
YvTa4ivARRcTIHynxyGIoiSQT/hYRT2yWvTw0j5hvBWWyigqb63vZlXxfHhBJQKfs25YVxrENYF6
qX+1wsTr/t6Y7BmheBUsSMLO5nggndknAt5qsx2951PNCXJI4BKxtnl+AdK2a0uOBBRz1YVuetXB
1P8uAqV3Oz3+NLLszFYfRH2Y2RlZDvDZt+7L3j0ixomH45HUXAQHe4c+ksn8DxRNhEOQ8T57yo+G
ETZx/PXKi4uuwr9LOzdcuvya6gTkYLvyepDQ3Ul4HaR8wPXkWoJglGG9SW1UaXhnFIpgi/lTXn5O
7u7sPBC5MAucrzWqG8cyhHWFBVaImMeyqH9zLF0WG8b20dtpYbJ8xIqfb1OJz7sg3cytKLeErwXI
SHhOrrpUz6NYZZtMztmaGBkk2JYEX80EsdjBuEhEUI/QZ1Umzm8Yv7H4pzVHWuIaLQp3bIlUHIk0
1+0y4ZWYKJ22qVaPFbpsfwlNZ0Oa5pzao0S0ENQpwF5tkldRcnH0fnCF7VkYrxPRQttGjcLguPM7
BeFytxqrKwcbd5SJP64bK0nuoR5tcg14zsrPVJzXZ1xPFHfHIpPE6/JA2C5lHBuGv3oMtUrdqykS
2c9OPqOKqctNI5QqGvnkSunBKzBaXxHLJIY/Fev5jmrHvOD3AuTxKCx+YMJgGk0JetiHKmad7AGE
CAHqJyTT4WC9LzPJkASumKNDLDhy8KxpaOsE8ieWFwOQjHPUqmK+tDT+FT34g3AX1MOKMIR16ZI4
kPaxW5ciPrY0lOrvyJPK6tuKpatB8TWrvC23uoF2rd23qQugWI4O9ltFnRal3NAG/BHGMHhdPCNO
fOPkighfMVbyR7DjxsioDFkAIfwfxq3RjBlxyw0jTIiWW197zWAZ/UoUYtnY/8M9Ipk+o90mxXzm
GUy47jmPfXI2uufKsSqPtZT2IlbwpfYE4Oo67hn4TH15OeeZyR1r/Y3Fk+iy9rsq1eRZUIK79l4r
4eOzoCnqJSsftKjA7XxwITtknZ1GHxCMuTmI03nL45hKZ66KqNPMWHz9Pw0GLars/EdHMU7Avt4P
BF9Aek0qRmWzzLbi6fzv80lAun3QSAXhzYzMQT192XdGX1oo/l/SyeC8pm8S2QxYhjyDH/DjuwZd
9NW9swAPpWEi3979ooYC/mm3HC3nide3nJ+PqCYD4+8vZl1Jt9Jaq1VsmZETUKElZWmzL2YHVgJg
AitL99LjC8kJrnnxVlJjfHMk+rASrD9SzKajVUqOdSXMrHIWRh8ZDAf/mB/aB3pyWCcbMzmnpP4f
kA7kp+/d7tgLLIL898oO/eWRf014P8HrwmfSOFj95+YiHYmG8Vw6C3wkJ2fKSTMpFGj0K4wXL1P8
kPuvz/jEnX/CIXn98hvWFUrxtXOckzSF1Urm2iMyRuuzbGXD2b45o39DvrA7shWRXI5ZRH0yo/sh
G+KLLWjZ8FywON+VNqetIyMuAlSf0qhgIGq09Px233OKPXwSs6HxaXajR+QNlMFccRbBSF8P+2tv
qNA+oUBWbE9yib7GulxzQShHX7jT2EjWi2cC/9fPOfEUaZrS0oBBYfdNcjlTQ6c8+P38hRmn8gRm
LL2Zari6ligUYgzhU4rQBoliCRi/xlSYT/oYN74/JOE0iVQlJkAe+5uby+77FEIQA/iIjb7/lokx
z+69UJNLhfEtk17LCw/NDqGJhEP4gw9UTsS+3zPqLarjHN2JWWjWvk8SgLxS2FTn6rR/OmslpJBn
BZbcQOVEd/VYmtUnhXcbCwU5z/Tdbfp3jjSbGwT2X71galOmLtF/W34fMV5XRlXoguMU++VQ5Ulq
XjSh/4YtBEJ5gArKY3f6oFjQ+iZcz/SZ3NLDeyHM8KK0pKThokV1HF28XkMXzMX2JTN5+1lXkRSf
w5yo/oVHZdrPe37NIfPZGDMepm/aY6dupQQ5YX/d9cQyxrjDGlgmavBCSw+tUGkWSxGVpk/TMmzh
n+wYEWbERjrofW0UzYwxVnp9GTof54e3cLvtbRJXKhzRiA2c7sA4xRhX4/uZNY2YMaXDyOd4FSSz
B4818hWKAEz+a8f8w8pwHHHUSR4fvDUviyUNlXauY3ZohEeFMFDq9GpsA9/Y7EKI4OoFRQ/WLQFB
chz/lvYkvQBEuWFu4QHB45Ar8lJ8HUAq7JC7eeRjLiPGu15upOSulFmkleJYF5oGlrNX2S7GCrdG
Sm5yToa9SVJSP9bnuFtAY3QEB5IQuDe0P1N97wJI8DXbIxMU3mijN5yW7hrBIKihciUyxnlsnbVj
AHKkTJCZM1mup1Q94TcL4yk+g2j5QFzCAKgKgkq/qMDZuJDzwVJoMieWNHHeS/LRKYDu1yU9xZLf
Cql1lnWfQpaqWVZO4di5frqoIBJqPWoQ/hFWf+v16Jm1Hvbzwbc9XryV8RKfH6pEeOOLUk98j8DL
e1g5Uot8Xh0so8SMhVtK7gXq9o2HFwF3ywo4w3OBgfDIvFUhxJISuYpBwyz20c5pvaz9IsDRGNCN
0EbnG/mhq0DKZwemVklOgAE52v3oJvZ+SvBvEty936C6bhxE4B8HsRjdio5tB8VUhAY2IIothq9M
omgJUFM63vBspIu4PA3QoElD84kTsjRga7jznRf8LM3975x0mfjpp5uk8JGkR+OgHty0nyZkeTNZ
8M12Rq29Cw7tEKR4Pw8/TZZNmu/BNMV4dFOGX1i4VKnjiz245x0E/Qg1b3UNAFDS7h6W7Ez0whM7
GwLlTCyOEJ15qxyPFw/Y2SDBh7qiq8FQLCwiCC4ZRkNj8QRrxHjcjyVlMUyq3sUY18Z+5buMowPg
qLYHoWY6X7mSdRCPvO3bmid+rf7lpI4An0t02qNnxljDprsfziGT9uD94m2oGV/1JAf88fLdSY9x
hRk3zrAyfGWOu5Lf8cmGJgbXLe2VkCxbfO/AtVOdNHNS5e64j6EOV/+gLhftAiasdK7ROJHnenin
rgy1Nuo5O2zqulXncuoVaAyPrYhYNBLFRH91WUJ4R2CwHXqqBkXwCbscW3vQw/j5kSZy5A2lD5L1
+9wQu1e6d719g7KTtqcqhLkLnxw4zjFAw73jEZLAi77Mv3+bXpKIv2eSy/7Dau+YcE3JUkPsnSbJ
m4XuY0UvuwLRvP6bMyelsh8iekNbkKHj9IlGLcOxu7QHfhZaPX0ZQPyUliamBrDr+0w9+VsMclqH
8R3DhkDf3/RDnkWq6DRsM+Z2ZfOoNugeL2E4gJohm/gJzNl3JUyZEjbcnz0bQO3VqGdDCPm4MRdL
wxi7g+xH47tfZ0O54oLFV7HDcDIN3R3SOWCjHveT8gpnda4KOrYFQZPAJX4MRZLt8YM+ib28MoVm
wb1Hmr0IKQ7h/Y1sC0ETJxiD9C6GlgWeDBfXn20AaCtDB72aJGpONPWYmI362swzQetuzmOKfWmG
miZtaRJKNcYCy9FLpicyBjkZSdDxlA/tlfaqVb1OSb9+OrDppnIEU2heoN8rO1L+YlyeEsXMzZ0P
XBTuSC5yg9luyvWVnb9Oj4HlYXDMv+9w1O8ktTtSwWf3Y0CmWVBVEHTrP83ui/6agm0xsY48EFv3
CpD0hwPqAEL1XVsuHO+qlgbobrEIJ5vsJ3kq0aRpgWME4Er8YQUMcAXcAUzH2JXhnuB3uBC/A3mt
ilTlPBDZeFW7QOeXxB8FKTFDucp2Wkts4hk55PppJ7nyduaxT3Bz+3W2zSBjFX6JfICmuW5WzTOe
in2/cIs44so6XpFoxlTdszCDhxMfGgj7WDvLssIXvZ3NTjfOk1cYYPNmOgHK7yZMPpPS5bahhns0
ynOG8XUG/1vZPmCFWzz01IzWMa8qHQOrfqNUZPAoAXB4bXZvGZBZwliKAf3OJkHMlCQwzdqsq1PW
Bjzbq0PJ1+IvMIjX7ast/8TQXOk+1AER2Ralv0OtQlvv72fPtKK8bBIA5RV8iGfDZ1dgGu1YBc+k
WMBoEydIxw7gvj3c7Os97v7AAc325j8oy8H7UZaGjszdUcLxtS7H0GGfJsy/T1S+ye+tVzvmYGoX
UzxX1FSq3yB7tM3Y0Ki4THvyMXFgFWPk5DXgKPlM9IE4rN3+eKo7FCQKXZZjzf3vF3dfmbugLfgf
q79N4COXx7WohHtQ7ugPXLArlUeSzMWE4mTHPqX34uX38kPZ1GNrxuEHck7+E5igDxm0pY3x0pgw
8aKYn13Q0+zvKZdQRjicsVDp1KqgG/Q/TNBkcYOmkuO05eO/hdHCFKevPK8DHLudqtThkxgsxJ88
Qm+fIZFEQGiTNANeKI7r4BUtj+Qq4CbbbCGUzhvqPupZtzWmx1tRIBLcsaWyqzEHXkLDf7/ilOtO
J7uFbZqsA2Ic998fhpd3PnIEDYppEEHFHgjnxAkRrpHyMBuI9lanqyDXXuxUc18Ea9fBqNT/4cpF
h55Me4MEtbCeLW881d++NN5d7lEGEom7aqnG8/TIW4tWi8LvVBhfKUfHGR3CXVFaYYeIZKk4Aunt
I1ubaLc7Z27J/jK1ZZWeKse6I8txMby9eeU20OnEIV3/fIjVCCg8DjVRzt6i/7Hunz05S/icD0CX
kWjVX7EXpqIhfRY56XBCbeUPjrSKqXGGmEaPsKs/ZBU6VlqGzBlRBCcCJ+bWrGZovfJ48Xo8AwIE
rrTan0YC5zlUmtgP5ic/3jO7fEK97UA0q2RuTCLScbe10F7yfHoui36qrmNx6rgrqpTW/VsGgk7e
RTrysUS4fIyZOQP5Ja/0Ga/qYoqdxspUgt7ev2DhIvrO51J+7yt3h/gA+cTLTgnkxA4CjKypgu/t
M3IX1DIkclsRMz12ef6usoETOdeVYMquwcwk4kiBzCtl0Qqw6tq0AK6BMPiRwSDeW8RSR/jPoNRg
ZDWGxuP+m1zeRGkXMe/dDqN/LYeIEGfZ6Gvoazeacbs6QcDoozhU7PTS/TN3AI5MnFs1S2hIntYm
ud+XtLye+Z9AVaeoVX8YOWBigc08jCE5tw3PDNnmH2agnPJpSnwLMBoqZeoXUyz6Fscl1uQ0wGJW
o0I+UqO87bMZc4qazE6byoBKSEnvlLBifXtVzchWszyCxOytVwhpDfIeuAjA7BJEJqE6gLfmEFJy
rJbC8C8aBoX6Nsa/Qp6/qR7IfdHa/QaHerB2ytazetBuW8mR2zr5wshDvgPIr9zGxrf2rNhdJJiF
yhmy8qLdWx+fvpnl5ND+OImv4ySta+kPU233OnrG8iZpOpYFCvbKbwu3MYpcJeTrywrm9cey2JFu
pF/WTC9JjTndGQEOcZ6tSYMhOibTy8a04cJlhgZdx5ubN/JA4/tYcbpQbelXXfyJHB3Cq81iLz8M
HRtvIdNWuFRfOyNuR8+eChTFfBnh0Vr3ShfBpYcFGYo6LoyLNj0HOsrIUEh/L6XVTyXFwcUyTYuF
sENAItOMXMGd/rkjRVFARGqDt3HLbvqX7QxmVjePjNUzYFzhfyzrussBIh4kRuE9nt7G+D1w2wSW
UWOLwftmxHUGNmD29K7H3M9mfRj3ug1QzZhjmDRCQ6coBY3SUCVwlWE2V2H0fc7kEHon0hUx7l0/
uYkbvK+T32/JUn8rrezScFyHmG0mT0A2EYo2wLmnDSEBW3MdPYUxll9J+v/kYwYkLCnXRDsm7D5m
gHsmtAxNg8MfZoasTDkt8GB+EXK2NMroYFUC6XTum1EByt1K/Al/mdKKL9nusOUds4EgF0hw2XA5
Hjz39DPdnxmZk+5a6f+G7OeBL2UN9q6uI1tPLrl9jZCNCg4SSL3/vW33/kXWkcP27gDUykikVlar
jmPgfJLLhha8oxjSU/g1ic6J7pIUbn69K7ObKxQXTfQ/eisDdaHCWZy6ziUXZxbj9mKGDE+4z+fE
fvd0DNCQJML3rgMUjvEnLadfEhlQ99UucnVfVVk13v3LEZP0ZdYiEJIxzAXOMsCV6Q4fB0d27Ava
b/i5cwVwviXa+cjqHzUIGRQ+if8We9tnT3cMjUJkMr2bHs55sJp84IyCvBZduxszcURMUvGXFhzK
d6s4B/b0oVomzfbyaBzGEvIUAsk2KcxP2Ro5uXHyIHPfXlINS8zS+sgPNA/FaoNIFsNU3JhfWXHn
wVlgk9r2n66v6pv+dlrnkR5LnyTqIyPxVTD2R3bqVX7Fp9x9lrIwhaosqV16xxwsXBTNE+/2ePXg
rbdlNoEWgpOIut4yGbx6X5aS55d3oJ0veeUK1PwTXZU06VgIze/h2D791MTFu1JVtYK7tNKk4ynj
puTsoCiQdNmTnTyN1HQl5Enr1aDPicTtQo2oMWvV8V4GAtS9yYIcsZLV4n9624Ko8/jn15Oyik0g
k9MMEV0KPBtRok8wx2/zmMqp3QVAGvUMqOsnXQTMPAHyJNYsinB8hCHLbCL6baOGBkI1FE4/SsKL
l22+6Gsnbtp7BElzmipZHTAM78jweo9jdNLlUeRVf4bZYyJJRWgI07u12CSlMRSZyFuyzBELpTCA
iuaqYZC6Hu/OpGMtEJZ0lqRHztLJTB96HNiCPWqkug6atfCYXlQxnIY6XyxCDSEOMYTPnQ158t9d
x5qdRsLWWTDWd7V6yXJYGo7Rm7Mc6E09YkTV7rl8k3yCVLLo3XjAH3dEbU9a97UZgtfmv94RmN6H
k0B4C9rC/0qn0PhWYKY5M9QV92S47xahO3G+dwEm27e6zOPzOIH6lIGWgqwnxK3DCp4VF3//OPm2
27SuhFZT4zmX14D1PcsfcvFL6XdXzc76qvuMg7hrDQ/cKce56GsN07kTodvpxdwZ5DxS9gQnoQXr
Qx2N5JN5vyJwkbi9ZzyByNi0Htw1Ef8VzG0P9NHWKjdvWse15PJijA+ItflxIhFHKHQBtYcBfbhu
PS0jD4djOfp8MJ466Q+3N0wjsZd1Q9nc5ylRwohrmoxGa5WF1wre7WSM0elEQ8P6ADNjTT3igwCo
cHmcoS70gG50Td5V4ihocrI+THyOXsKqlba+Sei45L7YxbFZZCCHpeYLAfsQJMSIudyvOu8aGQMS
ozPyklC7ZRUpmkLgIknTtFra24jFneRMETl1EvOBZPRySr+g8DH7dUIiPZURkgiZrOM2dyJaYklt
pREG3yteaR1DY0dsRfSAxVgp0x0/vTKDyTjac87Uaw5RzdqM2TQqv+gWTI1g42THkJWNqpJbytR6
4mlNv/KoEGHz9kKbouyHzBGK45T1PbGmYv6J260FS2qnYLE6Raskiqn5zDAyEgZjgnKVm+D3B6F7
83Bm5wH6QorbMWJ1acO23UuX9m45HVo0FlYakXDv8n7L0kIyIcCVY66nrVILLGDVXGt7dri4KMT5
37qoTg2IoVy/JXpZRdWayurf6PpbEKpp0ULkgnUTk5mX8ptCfz0Y6frU5F3Z3glfA05R5VRBG/T9
qZVYEfZ7+pLH65dsD+Bl2j+BS90z0Y1lHYV7s+8w2qhVcbLMSiFxgZwxzV0eQezp8iOBMqhdKEKS
qiAOukgnKXjW0ivQ0NWaiuIHu2Oz1NQeAlwvK+DkAPbOHdUnxNY6FmdhigSanvqfmjfVpQj2Ifrh
h/Wtkvn/nfBquM06QdDpqvKGmHoFZJgCjzmK5H0A4jHFxV1nPzUaC5w88EkTk+Ap6299rVFkbym4
28/GVg5kSOlDSJtR4/R207XKlGC4bDt/L+GOMPcD9y7ecCCLD41md5HKuWRvWKmy3O4PwgybrgqA
smLPKIzZ2f4Df0BmYlhDiAIBATqpNed+4BhEqUz/vkzZU5ZHEFaolDJlXJtocVoGltOSGZ6q/ukC
5/gnpG/AbCyTgL9cpccStyRmEu3yWmuVsXw1/l0QNidoNEKy1y9VA7KjPNSpzE/pzIV0bWM4cJ+L
srlDnH1csT3OF6sotv2Rs9u0UHrSYuyjb6bHG5AYbD91N7d7xtB3bsdOxOaT4XRwafwDJVfXO4VR
KliAFhu7vzpOnfTt2JaZ65Po/HVoODFIMZSmUtPDrd7+VVNFg/Q+SfbrDtJAWk9qECggQO2MKl+D
QnNQta8CBM1DzhfJPIsOorZGaztl3YqBHxx4ZHE4uXj4k7u2PygSyfbrw4xG6jJyJBUJzvaCFDaG
pdOa87ad8d+nDqDCuSAuZsc/fh4Rw0xoZoEEi0B9hfq0FCwxz9egG1yrxIm686osnVU6LoUgbJBP
sSnHRDA1NC5T4nrnqhmZcDR0fL45z2s1JPjWZGV9Zm0tkndHeDjyhPDSBVCThLbr8wwrx/lOnk5U
JsDY8epjM8Aq3LTlWYlHAuzpqSjUXrUDdlw1o9FTChtOEV/Lp/DcUgISmU6pUnQAnZD+dlEGmsH3
0zX++sFXH7F4KmNPWa0ZJL766DX4HREjHXx+qXQrxIuWd6Gze/2tvfyhgxLVc6ic4AZZGUtdqBeH
vwPvLQ9ROS4twMejzFBWH3zKjFtsNxK5r5LmYUzWH3AVmVddSiN5FFxWObjBAjTORr5iWQSpMYSL
ytFGmvYhttGIVQg7Fqu63OG6Vn/QiRe6X6lGEuio2HwcV/ceUiFiitCpV2O9hn7+uSXpGY3SbkAw
hMdgthViKbG30AC5cRh5wfjOogFfkWCTKjGIgp+X87A9RfhOc3ycXyL2xDZXCpCRdz8fiIcLjEoX
dr1Rg2x+p+7Oc++fPt+as3nQHmXs2iYilRNGOYDDu1U2UphUbcwOx700TaaMwFXqbpeiVmiJbxc3
qlBrEp7HQiLUZl4Q48Q44AbsGxPxRIsWaC7uhTWZZ8TLmfac2X4TD4bHs2xUxndaHnh6jJXH+VpQ
hxXR/MzlTf2NqioK1aBeOe/ABihbMGuQuGErSc5c9uQ8HxqnShnVozA6UZnjaOUQZ/R+Y65SQBF7
uy1xis80+wOO3G1YUeqwk6SwJGmxxT9xndKtg4r1Gs9sNNpSPCv8lKVy7W/UqcUKR+DncYueyZBo
EUqVFVNy09f1jscm6tclZuIO0VM7SprfmeD9zXxBwomaKMwcqJTsQN1GZkIp8R0j+ubsjZcVdd78
s3YDisbAI6OULta7ZvJu36LBQRIJzU/m1X0bdDXm/y7IyzZt5EaGNDm4ehBXu1dFcsEwdT0hAQaJ
yt0DV7+SxvNuDQzcAgx1l6qGZFRl2jj8b2TV17x+cSCDnUDHCb8/ETdaVtt91waAuST3z0++QBx2
XE/XJQgIPHMzhntMYVGDvv4tOvkssj2jvw9sAnNqzWEnZxD4Pca5xXxbXMSd5LG34Q11fvjr+9ZW
PBH+2VoY37LgsmIOfZF8L4foRsJnmpU/zdND/dKPbwds1q7UitSXnksrQMspAbN/dx8m0H3wgwxt
sMJ+BS5RVLAW5j3PF9vBAMR9fyYFfrBiX5fOV94Jv8cPTMtp25pgtONzZmMsz67yyZAwzjb3Llfg
MQG41Fb6uuxzk13HaZ33ZzHvfigw78Z7lSydqWUJ1hoG7rqDiZnTiC3OfG7Lkw9ZIY99SGMRA8fA
eI8fGRbdjoYmqsBHC1ODStuc/vk3jV+VL8sAQ4TU5vM5Oj0OeHv6gbMDWDgcpoynMcwONMHGUVAV
rRZszIsLwKBiS1HurIHDREJ477wkouTbkqFeG1YluPedcoEEbWxHTnNDEDFkhTxIF2JDNlQ3UKnL
f+1Qh3zodEw1kxHm+iB6CEbH38+0GHaEwaVhwOPR2nL6AZyKluTUnEFlIfWLWHz/aGjBF50TSjn5
N4aIMycTKtI9nyEtzyIZS2xIwkHk05fYR4MygV++DwEEvbYWPqnQjKFg4ihLV24Q5UVNILF0Da66
8GwPw8+So2E76ocUR4m4SzTKYbRmlwyVvIEYWo8ucvL8v8s9Uw8VgfkqvK9Rm/FI2eA1Z872yjjP
IBEku4Ih7PZvMP7WyrV/2Frsb3tJ4PZLWyNNg8K+ccxKXA4B0mils0MiJN44zdBWVjPFg7aoktc8
kch/0yvNIZJiEzow6UC9K9bHy4CjAecgerolxstcciHONgCVUOjHhsjXMWP1gKACTmAk/ecuKtqq
2B7lzRr1TJN3QadabRUT0zcR1b0BRqUr1HIra8N2aKMl96TG8F3ReTmLes20Ohnezuo0E0z4z3fw
F1/1iCbVOtXc8joCzGkEVpg6l3IWh+jlqz0nkP5f4nrGk8de9N4rvQPO2xIxFCCoJCAm9ezNSt8H
WariQr02ebr/HXiV71cy9ZFiQnfvlPCQQ3261Aq2oWafwA2UDufszaMsD5Zr6XQjA0g5OUX5aNYn
EgnfSj7CeNuRXBuCTGkw73mp7iksijvdSXES+AZCjmGGYaw0i/VipUYd+4vBNZHvKrYxV6JIZpgE
ZCselBeM7vUrotUVVAiuqid6dYIXBcSWyhhKe355uTzKiT20k54nBjxZjhsIMF0JkGyxRhng39Fb
4rNEYCMcuArcBeOykrdaYMjCeRVrVwGd5hQzKiK29ieIjOvwYJ5TZVY5csgx+aiNPyChlGAJw9k4
wTD10cu7Oo/z2CWnDwzKGCqL3chvSskjrBlEwYdAjIjnJKTWqMKxF1hMSbcx19l1K0jolEm0AhEU
pQiC/XNJIYx5insfqk2q4ilupHsJYqp0ufH2XLjL9ZyGe24JhAv3m+8zjSDUXUm0SErAHYHokKK/
zdKdXEYQpzYFXys2WqIFRrYernZZJwDOityccofiwNC00XUR1Z2uGb8bghDKJmNiPNEbzfIp269o
1UsohhpXE3FOqjlXdtqAmaBIsivKWARFaZLcxF0qLwdebJvu6Z2JfSCK6eG5tZlC6Rkac+KAKKJv
ouqNlpZejAs8hkJ1ZYmw6BtGqiUgZDjHwzRRUhaEKNWB97yxKDND24xG8yfYoFdshjWVysi8SwqF
KjOoVveaWPK6HZCJujJktgIPqH9BwDLPVaAAFM321nGcvPDwxSXUL3beauhrsmx3lP/FEjmJ+nUV
bSs+/g3SnBszL9q8Yp4nIrfNvvXZeGFqcyFlCGyAWyBc/yLYya32E+sPy9aRHVWAsDUHIymrQKWt
9r1Ti9GWKMjGpjFkIiCFFeZu/gvX8B4GkyuFbrdl/1DxvarlJX13D8a23lM7A+UxaHiA+N4qGqM2
6nmaAdiUIJKU8qGYEC8Fuw7zRgmV63kWua0on7pbuos/Sg4L3ODFi9BytMJq4WGabttTcaM1+SL3
LdVQak1jkHP1oLIoZaNNuvZh4KIOXHbdmSyto/p488NMenY5ciDDDDDTeHRZvRTUFwilh7VSIxVQ
JmJXMIm4sxz+dxwHwU4a2AdOhMj6Fiv3qiP6I4guNaVaA+HJz0IExRtUEC8crb0heUEmjzOqPY62
k+HrnGDnLGySceB0bb9FCwOwfYkt+532MX/XRZqOH54iK+ytL+VXuHsMFxOqar9jgBNNaRf30wen
5dP5kEAxxhl9cxcQE0fNziaqXNuuT98QfrWZoJ7UJC+woW8kHfz+uPOLzT6tN/G50LRxces7rQxN
18HcN5WTY6iem3MdMcQpWuJnjWtu4lTLaLl22aExUWyu0BT9RosjTsOM6gcpQrmsMyZD2jeyby2+
UVEeTOSXUTsVLXTWzc1Sa2Ja6567DxlWr3vag1pnZsYlfSn217dvXm5drcykc/iwa8oNrEAm8sM5
X6m8Ee0mh0gBafRXfcaeg14k7r0wBFJvOA7eRAZHkXUa5vODRv/pANBUhjTAmbTujtyIMtJFUSt+
d1Mlfv/gkgZGSef5xEafQFenzdAWuI83uyYpLVOONDmsbh2EJOjOXe3a3eSdNxFERt3QGrWoyVsu
IuyTxmSAnVyGiLhNJiWcCGAo2ZKtGOuFHmHX/4AeR5Xq8wCXDO+7UqZy4/cFJUV8BXrernrjiB4/
I7OpOKFSuhN0IE2igGuoGMfiQvBBGuphiQJ5qiV2Co/trDx7PhMWGA+A0I2/XzsTD85m39E0UAQF
9I3jj+EgMS1KvTAN0+yjF1TjMIGNhP7D6Gwd254zXu1uOXBpbKdZVFfWkoK4BIsF5nQS1I9BdlFh
vXCZ/isZxOKEU/O/h4QqOwLgEI4Y1e7JGOe6u1hDzv7pHrMsa3jp2kJhQM6mJUVt5rFxuHxc4+kM
juYOWjDGWKDbLOlQGcmjEdOq+7lI0S0ZTWPaziEMiS/hE1dVNDVRiAo9fJzbQDxdNHVmMRAvpSKB
Q1sQpi4XbRHHP+suy4tdBLHxsa9BHIst1CAo2wNa4qUjIpiHEv/aH50Gk+tmslgklBn+HaEMh3SZ
u+0LE6H6pDb/+Y5/Cmr+emwmCv0Exf5/mbDoW79gufFKNe0mPL0qyRX2FXZGYUSpUBWbnKf6zMaO
NbPMoS7cDNasM02JIDTmEl1WKIKBAtxRX+5m/l8hbg5FsHK5KtswWP8QkN29zLOfvBopb9i0g3np
Y1cxTvFmueohzvgxD3bFIj/OPqw8MHIgSHZCfIanvPmJjguNn2Bm13Bl2+Logbrt3B4zV34dqFH0
ji0pX/CtGCpdWD93ZODijkx0w4gU2StmoxtSfKkeBcKGrQ1T4a+9OOYBLNEVPan2KABxFCJvQByL
beKEuBfLTF7iccUzUH9jaYWuIvsvCNcgAopx4JqtbpJ0JOX0xcxjBrk4Bs64mbbEsGoNzXBaAoQb
xNoM+ze+RyAL9A/zsR1VGA7t5/CYyxuAUf+Z5Juf1Ma8WZ41mcb0LaXThXY2GuDMZC1CZVA5NNfi
Q+Z74RZCoLkW8nfuh/FOYmJXTbIfgDAO00/qoj6CSOJxzjIS/baDP7TpAmaUNrFHDVOD2kVQxDpA
GOSwew9GfMsvnfWfLMzLetjwi7khtCctNMcP/xGrg102D0Mjh3QMrO88AsPXUFtUJaYtEeF+pwSm
GCLUp9mEz3lZKjKrAFTajv+qj2vi03imW/tlGqSCAxWxTKRqBBbIQzVfZey/lQMkMCysZf9ZieCh
vzBvy7Mbhx8Qf+oIpyjXog+jKrr0xVf9Q8nqlXP2Kbf17XJMy0MgoFHelxO45IffnL7XfWY0tkC2
qKjOFwOhl52cmaTW2ibnhRO66YxCGwwcpBZcQNDxvjQuawyj/E7JXy182Cfr7zT1gQgfQjtHWWf4
VRSt6sYyJ0BJ1CvwCkwZ7nGOT0Go1gharqTQq2YMBuSiGZ/2YDYbYFY2EmULVunLvs+fGmScdE4w
JEPSdXnjS2wqyvTV/CuwJkDztZvA1YCbTUBqqdyO12/knSCz8L2nuneM9PT7/FM9j/A/kiVfblfY
lJfNCqV6vZR+zVFVNCv9azAQWawisLu22gmE3rWaX4X5pmL84jXqeesr6+xPTFy6np0BazDDFmfw
RKRlUJ1nI2dObAMeo4CFrCH/icunTe3CLX9P1pEagyBsdF6ATugF0fiHisxumxIzRqn4Di7ofyXb
6dOE8rexA8wpyYak3/qqn/AIG1aXaeUyXXGbtR/6x3lX9oV/GkeLIMokF0E4cRvJlOyWsTfrPy0j
aoluf381ruNVYUQYJTEy1GgM614neyFjwknkO4jJHBeQdkaoytkPGHoF3hyUiOIHsCizJMlCRj8Y
u8ZwOYrOP4Nhu7lqrpCf7jfpOUHBDy5NMrrv6mUGqqWo6UoqkSmRvVQKw6NW1871heW52I+R9qPd
7r8RKBXCas7mYMj7sBIQcfYW/BL9BpI3UxMzylUX97A8YeWM4elD5JpPisfTEbdAo62rAzP6L9cg
XY6ZROw3fmYCf6awCftGfRpDpxSyaKMdQ/ZtU8CzSQuF1f0opRqnn3Vkbvn0uHHuMVa6FsJ7uZHP
Fh6soDnTKJ84ff5e3MK9n0IyFjeWBb29XPdvo6fYJGvYJlviD1JHDkU9l2KMMgh+RU03KdCm05Qm
D12Fvbt9IHqxwNQymTqDPMI0H1i3EhqzJaVSW1EZZ31e1wmE/sFAf5aokmbEMmhEW6XfrP452ho+
toLFaxxzckVhlZGwke+ljbCtlfNmivF48stoC5XOd8mBXLhF6maozzvn9ERAHwYkIgfsy4L7Bqu5
oBT1FVZHCYdLICV23vCfb3K+MFc+nBOmolpTUpsRUOgPZp6JwsJJlbmlnLnVBc0c+4HNd84bOnGn
OZ1cLKsXIqBcJNpciwy2Kf+0DgYBo3rpTWgA/JpcAwZnj+nJnpaDcm1ppDXQPXn20C0C+NFO9rV3
B9/7CuA9IVbTvjXua3ljsksc8OAMWsGNdX5hSVe2Iz6wAOrMbjSc4R9EU4DBK3hT7jBxoOjqECyi
dcTQP3XYYmtlk9GxvMLoxb/nBjwsjZiIYFb4cOwjTlRPOrhQFIop+iCjS/Lp2ESAprmQYE4mc5wb
O9BjMUX5Er2nE9TDNi+HS6V9LjnJy4Pw3VLS4E8ljq3DC0oLymkml7aEaZZYEhQHeWisGNNv4SjY
vP0WmKOg1aKp+GNII8FqpULnmmfoSYjwEbCiMhodrZmh6rzWMTD5pQtRP6sbSTxaGuIXSsTMwzLQ
MzsVzktPXyr06f3v4/NDnpx4gz5aSopghyUP9RH1V9FoJzztxiH2zEGYqrDT5fArNxCOPxiFZlQ6
q4vrhCwoa1DdJ/CqxudcYubmup+peGE/y8vg9gK/7lCZ+vgWDBV+l485Na0N83NDok5LDcadEU3S
YwjB0Wt5j1tZa3lIy1UZQTfLvYk/3wlY6GWIjnEY1gUnOT4ACdE1oGYTVQ72M++4/y9k0HMEU5TK
FD2WABCNG6LBHR+qTcE59H5iyPSuRvGOZxUlTR5uslvK1uQu+p94T3CdWhn+ayX/+5a/LYqjxDnP
t/zTxW/vjGiWl4O2kBvyPb4Vx6IBd3d5dX/Aq6wLadMq7t3QkgI/0wOVsu47QpYy93JQqtHtyjlG
wAUg26utPcqH/j4DK/QsUf1LLo3nVfJTbopnP5gQ6fmPOziQO2M2IWASMHXR09Mt9V0gq5WSnVa7
O0klNvOLCfBuU68NTm2DACd48hKwM3CDTNreziwyQJHG+stH9TB68dmXzSf75gjT7c2OXnCsQWsJ
KQukjXO1iyitefMgbpJCAvE7aXJNgzH0UxVGw3Hhm033rEBCb2HOIHGMKDzzrek/mz8OhqQcGwCx
kK9pAwD2qlJ+gqHwihxFimBErV4xhSaKZJOQya1xlnydgZnq5r7vxdW45Lt1l84jA9Pe1VubgAy5
ionWdjx4nSvaGV+CVwrf5mSKx/BTniu2ZvdT+G+VAva3BDl/6JFV8EgFA0Y7DTR986pXO7YYeM4X
w8LCVJQGu82XGHhsCjLdepHplnK7VvBzQBLMTiE8K5AWsf3ph0BQk7JcriO0PToDQGe2Fuj1xT8n
5GnAA+yL9psN2n/BJwANwzhCuhrEKc+EfjPAkc/j1SZGvPeVVrivH0FSCAqK4YwkR6KVN+/dhDUb
rPOqkq8s+mfHhJPIEhY2/Zir3+GMBrhNsN9VGNwqSA6MIsaoa5R110te6VyFt5O8xHLZ1H9Su7Q4
hfKmyjFxx6yAyBmN3KkgU3iPfIzswELCJIwAONBgXErLYNE7y6DYYKJH8EdSAhr8wUCYWfhHhfhf
IXXXV9bCN9+wyNH277d230lWQQ0JygqtjVQpOu8bx7G8isaQ2JTMyjfitCWI4KUvEf4K6Uhhvmy5
lgNigdsOr/Sd58qN5HvJpaQoa3sp0kdjUPX9KSUbsNI8FfaYFXNgHpur0oO6opeArzYrwA0EK5Ea
xMEbwPM+kKYZ0i6NTJB4vdl+e3DVp5mfL6AuQ7BmKAGmpYGAuGJbbKdtBnGx2lR6qLfhPWbs0lgY
q9jKTJcxd80dDBS6dDIvnho8zurFUlyfHbo4k90Q8wKm/1T7EkzckWiZa04hp+4GVQ2wDYAiI85J
LMkdIEnSqjpJsIBTFCxkPE7bM80lMAZF6xS04QF3ul+nmfwJwC7RkXi9wQHE1Sqy7qidYegb9HkI
3//Pzwh1g3XHfMiJdGRuoMW/5fQl+ztJ1MxJstKV5S1f8pNN1h4qThrFmg46dqJv9dMUf+u/wihv
TyXbm+NHEL6Y6lSPKWwCjW7bRfW2HDHk9aeQusdWdnGMZPRhqwOoXYRdEsJ7SmICRxAr/YsKqPd8
Uxe8XW/sjRZPz5PlfJXUTaumHVYTm/g2jdtz2t+7zPKCU7iJKlRfFRKFqVl0H1hEtSowuZcwJLYc
pnE+KMe/Kjra5Hspgr/PJAg/Uj+pUk3Q7xt7rqstxpwfAOvBMs5H3O+VdXT+Qy7SeKpl4m5aOGxH
jo5I9XRbceB1Ozd8wxlUG+7EnkojNGO5jBma97YpanTDiEVzDxG6fgYptG5Cy5lzoKBjw2TrHkZy
3UlXvxU0IhpiQZ7cCiCm/rBWJUsb92zy9llNjpE0fq3WbtLEdJ3YG4CcY0eEuI18DdkOLW/nXCIK
BzTbGgtLDqmitBblnSNaEo/7+E+e3ndRjy6FyLJb7pUN6UFWr2I1L1RGkeGv+3S5LG3t0jQ3ueuO
oDurAi54u9TEJw3zC/q2tzNfdar5zU4vhnnABs/cuz/P2Q5YaDpQlUkCwyHXYWhAflDaxipPJdsu
rfcjUPkiRoOO0tITnwO3IvECmcMKS5Lj1/BephH3anEzUohZVoHVK9Z4efOowziF9UNyoTpV70up
WqJ25LHKIl6QZ6QwpVNIGJqxzhRx/eFDvYKFlmq4lmV+XXeIv6sdF0FkEvlEYUgLUMikJU1LtE5k
CT/tjCp3yuBdWQc2gRbtGVu0kBdSnkM+KPOZtEsp4swcqAdbSTaKjvI2a2TGJYiCuE3M0ed7kDzk
6z/CbYtdwdYfLy26WaVP5w0cOQ4RA0LxkWQYIQkxsl4pMdPFZARPOB+/YjPdFTdkrD6gztESm9Cm
HFuG+rtQf0if2rF3one6kckRFWrTl4xLQERyeXGbXTYwdyUITFjFckWJk62Qs/zI8zHt454TK8tO
9XsPRIkhbeLQGlXNDvLqtniAqKN5mKwaOnyoXD1zaNSDn6EnIEo1P5ZmewZ/SQlhIA5rth4eXD7d
L5lhNhmOw/uf9+mMRxIjkgBGuE0zPiPzDlJWnFCoh3aEerxgEHt5b3nE9Wlci6IkSN9m+krod3Nr
SyFnVLuutwCBkQAwzWwj6OGF6BXORZPAa6BuLwH1bf+a+T9IhfJG6yURyqTZm21pj/3li+RG5XCl
eZF7jXl/s9VsepRqH+IDU6BOi07qBxHZfZcl93QLeW+2/ovQ62SsYoCxMJHcgJxjyEPLFy8FSdDB
E5dVFrH2ke+ceIhSmYSAOD+st9Tx22zGnSK75Wj76AmtLNKiNByHcrt7G2fnYQ5+D+xJNTvBt215
phI32pz65wu/F8+7iN5ZzJNJYt2Q4hbQpcblRvyiGQB6umkxcGmgMxIlZiWRIzl9A8bLJmOgRoNV
LYiIzDGiMKM4rRyQrcaTnLTd56QHm6PUJD483xq3qVBqD9pJ5luRmqnROQL6KbcAznF2jV7WgEje
pri6Sgs+i5PL0BbUKYbhvr/lnqg8th6Hqwr0bZrUellpHrFBn0AWAOZ8q/AdJCrhu2P0yuzW663V
/T0pD1w6oOyU3y5WXbVnXmot2svNAqg2UFj8sfqmQ6PcIdy9eMvQSvsGyCFpafxHXUJiBlmU1g0/
CHL2UnwYngz7oQvcIxod/5d1dZ8gizfj/hyBWZWpH3SYyyJN52q0uCJii8aQMFsuIP2CNaDsRPNA
gr/0RL/ftmT0k4QoveXs/evfejndIaF8qB77PwAsa89EfzMb3Ae6wHk/BDsYClbT51Ye11/+iMDe
ZDkXbraEJFTclX3o+V7FA64rmlZF7D57E7LMb6sSDIPZ900gWmMXJfncuKRR4damSuKmi3z99saT
x7r938dZ4+iOMB+g18Fa7i21gTx36alQk2mfEg1WijsdBMi7GnTm1QrZ729ojYfoQ8FLiiBwDniS
QRAZybPNEf66fAGhXmIGuTnX4pugNC1jYfLl14ZyI9h616Xtuzi09+/TMrXhT2BS+8O9TlyWjMr5
ei382EsjvgwLptVeLQbQ/vlsCrnQUrbEYSWThI/trVazaKGvnXu1xodP0JCHwQII/wRs6TxoBBol
UEl4mY0418yyveIUYCWqa+FxP6YBF672RoewI44gDVa/aY9b5dmuCvmXTxXCi098NMJ7PiyzNGXM
jojVvMfKyzrN5RdouyI1YpWooV9H8u6c5zgTckic4qVlXRNfD23AcHot7j8OQUISn9HNqLrrSD2S
ipNko/qJmal1B4xGJaanphp1fCPPSaLYSx5v49hiYp0SZRLDCcd7fuS1nYceSO0m7ov8eb4pCHVu
yx3xl3bXR9GSvzFHHk2UaxO67UxVhq1ozrdfUEvvFqn31s9Gv+CJmMedrabJO1oo/Plk7tSJ54YT
0vOlrkBQwgycC4v4BnddmU9eSL033cLfS2Oxl6rLUtpuAyvd4W2iCVN+Rxcx9kRv123YswZ90To/
GOome5HLx+pYkKvOksUD1x6l9Yb12Eco3tYPt7vBHtv9zFEbHi59UrCW2Gzr8+XeRsaitZ6ITyo0
s/+BpuhqqcqTG2YK+MV6eMRyjC36g48MJhfs5CmwPeZkLG7w0g9WwmTlrD6fQ+QG61AURDnyCMlL
JCJmjJ6IEtUdKh5xN9sUIGArlPB/nol0EV3EoyoZSXh3GSr+PEZmePxiVuAWSoSGTkKCwoQpFjfy
12qtFwSPUlTPcppr3QQejZZmCzNOb5byGBZ4gX8rq8ZX35qUc+lqnqpXRzKFzdiRHHWqUwhQY0n6
51L+CXhqP8AVi97XIg59HG5Gkvy9OgXC1MDiByyrr7Uno5vIOrNpQ7z8IsIhtVezeFdrMC+Vii3U
hfBp8gVdiBM2T+QS4yQuOPIIEZqQBSGZ9xhXSB06IUnls84nv/PZkupoYLLcRyYNnAaaLj1xxC/R
yz/Qlk2n5KaXShlXtdOZmm72VJwKCGRkIEccDNkmXNxukkhhY2fWLHUSHL1seca8o6XspKGn4hqZ
CGPBYHjsYebkkTidnhIzedzCDC4S+UKY3WxhTGTHKzxRuL2gSocUjnvUeISosOstRWxjKa5CuvHC
biWbNEbhMI4Tst5aXrHrurBogzMZIVNduynPSyOuQgY0WkdkHZzwMKkXyPEPmCki+f9dKsbvlpQ+
KSK8Kk1bYpQy17xY4iuDuu8GBPy8qkzJwqZgRos7gIw0LfiIFfURPL6c7q/IRmWFVBYXisvYs/a1
5umoq3bfoFQ3WICL8DSuLBIBmZFZPV6yo1aHxRMNTg6zWMFy0TSJTw8deijq6iJ5cpOt6DmgVjWY
p5IRVLU4zlCepzvkLYXuG2X+/I/MmRpL8N9kIzt/PuxPKAgDBkxYEvH0DjQKGjDJLmmcNt4Sd2Pt
Sr7p4yJMugubOQ4OS8e2cIKNDhEq+G6K6MsvQ2EkfpoowkCA7CRFKAe+Wthv2I6OUQ3ibKpNJySk
vUj+3WQntUsljvFQGu6Qbf9yCznMcHIKjz6YYV6Wi1jMqvZQ9vqdrJnNkEKwJ7j271a/DSkxrLVU
1sV9JLtTOMVZSOCmjLFLyT0Tz2gMr7y9HeEpY/menjecpUxyCbQi4419b/Ay1RqFOkLWH9/tGwMt
SdgG6fDx6n3r8RbU+GjbmDGXCyHsghfDfy04uVL/7W98U62mvNizV0wUnnq0Seo4uJMYrjD71nZw
Fqyn7BCT2vMKmeQxH1FaldFZA4uKKfQf3xnl2mJJQ6U7Ch11L0JtjjW6aQjBXQQzdgN+2IIFjdpF
8xpJlxM0eKGIZBoNW2H95UEnZJjz9w/3TFJycbBXHH5sr0YDoO8G3Fi67uHH2e14ckcK0iP3riHl
Nzm5aZEmFAcYZBVlyFPxQUuG34KnbhO8317zTh6wZNiIWZMnp7G6AnfJA0flBVefYAwrPbFieD+m
zXeXooJPsDWBWk7WIrsErBVsv/g6udnpMo+StG/Vo2rsr6U+wYiYSsAqwc9uNz2B5R48zHTI4IJl
YmIeO09u8znzblUC+WsR+Pkbjeef0Tb7YbcnW28TCXJJp/3nisXSgAQ+yH4NGbKegXXDZeZoefeT
oidHiYv+2AzUKjpzMXGI2hdEWqVj7RlJ7gKFyC0l5aQl5wFL9V2j2uYeQ3oLnANQJ+gx0SonTqwJ
kwac22n1OlwCckmrTJ4G/nFGkZRxfsPuiGQbophHNOVyk/+JVPKIBqdB0nFMKfTXed3daDknkysY
Mtd0tLceMI77JYukQMCGKoldeQq2axgJcZ4GWWZ4qdNcqfWrpY/UjDaZx2W/w1quWLU78tet5M0t
2xIuIA6drjz4m7OYQPd9Kw8TDAbaybowFbQjKQfFgQ55PYiLy2cB9xyNte7eVDJ1mZc4udX7NSuI
fYpbL/8+eSErB/s/jh99YYc1sQID8RMym97+htNcQ7TCc9ZromW9Riv5gCkDpnAqLlm4NL1a7pl9
bbNDsfBaE6xrbLJ7UD3NqZTNgGfUrWw9cHLSHrKijg82YOkIyylhxGRar+0a0CxZ1iNdUhRtb2JH
SgXwFwzCwe9YzNuavhI9g8bz9IKU/qfCmahHVCuXOxQdyMpSU8lQYReo8RQ66Rp1ByYqLSk6/lzb
zm2wHqAcCFeF3q8Mx/sjO8848CsbanwPmuGPGWhRymYNTPKIyIbEHeXFOTmmuJIrw0fPx2vNvoPK
whsY7HBEgdCjkem8EBXHhI4Oo8dtrdJFCmM/I/eqe1eXcZFNQFwUWZ4Pi8TnRIm6iZ2bYbpPeL5k
ineK5Kuc3At/JNfml33d/DSdw9cI1u8qvvcZWLsqswR4/+3meHTsHclwEi2M9Ye/9hhkz75cvgQm
svkv/1rYxZFb7JC4LUObcOCmTrKaqXtWmSiR0T/VxI7Z/uvTgTy4NZOvhub2A0dey0PJL5fza0vC
32PaZokSllFdHMPtNg7dtGwMtiBfP5udBJuu51nA3zvw1WejoX7f/u8yL16u7TmnbaKXIYqE+IO+
ZINi51vKxp7sdBj5oYK1IQFjPliEZWzwRMwtxZ3uKqHzZQ1p5r7cThNTXcAzCqakU4y2o3yOr2xw
JIiVkdrXJD2z66USMWzXi07bk/yaDbbwWdAfBo3Jud+ZF6/EY8O3L8IK9nHLDgdiH2BQXp//ksAk
7lpqdpG97m9r1fG2Ywoo7vFUwKZuJql448KpxL+LMcJEkYqqCzi7c82TYTjjdFCvcb2xXVearxdL
bBH3/9oV+ONSWgLgLaFcJcco5fUTg5cAZy3fn1G0ctzSrWvO4FmynLm7uhr1aDH998FDT5MVsqf4
viDK8HEilfi/zR1af/UJa+AkpBFFBFn/pwtzjKwhH+fsR/JZzGMUE+DrBOVD2dET0bHjFuRMkaw7
I2m3PXymEQI4QtwOzOqO0nBWM8wkbu8+FEAXATlV8uNbpK2tyUA2VZUgqcGwFl2NFr7s3Odf+5Tv
t79453Uxt2M+GZ87un+DYbmz5S137i6E4EMlsA8vhTPyCKfT3RSOKGaCC0AjKwOQac2A/HqOUY9f
oTZfp6isY8NTcvTnl03nZyNHEoK7cEja3D4qdZVClL342xW9vCdKG7VL15m1F6OBMB/nISxltJ6d
8nYVV18V2Gjte7iG+cYhAKvgpqyTR+85dQr9ZIxAfpKiUl8SCku8eECiA9YtSpSQYtSbUuVx8xCf
qpk7jkJ363F72zNsCZsZUggLHTJ/JlmIfV33SJ9276nbrKQMjB3fohRaECaz3O/fYtz9rvEiTUNZ
DUSYp4r6WMc0OyqcmJ9BsAfIyCp8bUCxsiHm4VIEnReJ7a1Xt4Li7dw50e9MQrb0aHssrANIRE4C
sJaMKocuMTm0D+9czaq5BPGZxG1clC1fHLSqbiTGZdJO84DoTHTJ57MGfVWRHQnEPxCX6tgleQP0
AjnLXhhSbvgRPYlD3knWMIKsTskorTB9AwbgztTvgfYErS2U9GiW65sEDerUa+vhO34dvOlByA6q
lnhjCSiqz2KNiuVMz4BeayiZyaFDk4Y5wKUlMssI+xS1tcoECDqcnfdy9g7w9l2KToN3BbI6zqNZ
MzQX4FoDG30ANDiOwj4FntgUnqisx2vdvr8m8kh9Irx/t+7AQYP1Lq6IQBUD4PlfnEBP7313EcJD
vb2j7XQ2sYWEL4BMKqUt1tA94uQbCQwPUGpwRvyzS/j0rA21JJkdW9cUqiVsEhrCJ5A0dapbr0I1
aRm/Oaj98tiefgfRtEdflEKrfTwJHr9kdKA6MA6eMGpJijwOYEUJwv4dZLXDr51UM7VKw07Di95B
69AEd0es1u5xREG9x9LO50oHPvdxjlfuaCgN4cs8jW7ku1QiuMEsvP1xopmQK9UTXAFAkh7EVdbQ
XuhR7P6VA/CXu9IE6wV4YoXaseDnNc+C4DwdctAElzNnS2diUR/OM0PSFUo+KGpWPdevFCMtvi6Y
T84GesnJevNXCNSapyuhFOtUREqBQ85dkZsdOBMEPLu093MsX9YxrEadjFW7AT1ARtufMX6E/HCC
SKHWmaQOepRYSsFdjqPAmDwh+fdTjIP8sOMIsi+iODEUhcqbbaFcP0XJMa9XP5VuinabxxyPbBIP
WRzKLpPwxu9HCXq/xatyZLxjYeJSGoiHG/f/xMd0jKtmMbCELzX/l9qISyEsR+fApZODeBeMGra/
DNU423koF5IlMWOy8aiP8I1bQ5qQ/gO8TKtTq6un3bxcasmsWc6OH2Dq+6dgEjS7dg7fKuKU3R07
pQyit+Vxu5hPAAxDMEarP5g4uLgjQc/0lOJ1WiX41HdTGvUIliDPAkHBYgAsQH+CgxBioC7wIE/O
aDTD4fMY3y3DsEst2z6re6/duNb2uDVDHpvWosswmEDD2hpWamDunBMqe9JDp5bDzsz4Bx+dKMHi
lh1rzlOk8AsBalsdpYDxmrUbGPqsFaQeBKdBxSN27zOZJ2U6vxNx/2ieUivfAApc020a6SwVp6Yp
lYEJt78OxRo+ajHNpxPDq59XbdLIYn74YcXV2I65XWYyxwArO5GOJoNHrTSk7Ke9/IefrzBAq3MT
Tc1Rnj0T6p0b0tVbe1dSd2TARAnI3o4QlBr2jnSO3qsUq3XGZCyAM7JdYC6PYOLBqbmtQ7SDaNKP
GeW/m0o4B8Q8vdG8tG+6UjpgyANusfY8DU+f3BjI3yILoGufJ6YpM2tmhHU74feBREgJpVEYcMR6
rUASmqjUK3FrNglIvoveqkzitiK87sDJwt+WX18/7pa007Y2nAstMQ+7kciThCedxTOSWPcxKgGN
weWUkwvTUoF6LTcUSDCtR/CVT8NABTddL6rBUd9cpTCKCstCi+Ymixmr7WUz04y5SsQxGgyGQ4LN
6lryRCf2Re7dTsXFDEeUgfTsQxfNToGQhNrJc+QNgqkShAOjFCN6NnE4pb5UpnUJUWOvcf5p2dcd
NDYE2jF4hh7eZWhcqGmB6BAfATuDQqfszu5oJEsIC0fGB4rJ4j9fho7dE4nRrE/OL6WZ58r3FhwW
B3qZH1qZNqZA6cAfYMq9xfPHsAEatO0uY62QaQXQ//vzCknlf4yzGoZRoTbx6H+5Gr7T0ajJWdw4
cQ/yGhY94fqN0cfynxYU5CwzUejv8E3zinwJexf3yJgPweylvXYTcZ1IcNDWwfOcF7C8yW8/80Ck
aO5rpIZawHcgMBqETa5hj/EQNrhdO1pdCnQldZLww7UHfwOUVuj3dH2CWVUDy55a0O1Kg/p+MR2q
wQxUF7JeEajw+bKaKWga8E3K/GtMHWUFg4HBbqdWwLjIZ8c8VvauC80D9Lfig++5I08t9yxFY0sL
5w/kxAL2Pq1sWcgWB0KEiJ6rZoUJY0YYAQukCV06kT7aMjNE/xpbmevOqh9oSnUKBQaMP+ZsfuOo
qsIBQg9ONCD/qdQK0N9twkSA4jgKjT+f6tBOywr8LOODc30xH3b6Np4LO4BItWtodGcrcXJEVxkd
WAVfmMF4+NhechMJcUnLNFxWPLG1VHCAI/rAHgAMLYf7on0pBvg0F1a0VsywG5TdJJEBncZA6yyv
LSemG/s9EwxhePiulMT+CUk/QiBnlKabSn9Pb2AxatdaD5Hz0fSd3D9TSxF2nc8rF5WmfGvh4OGA
HIUlh0Ka3h9bWb+1qq6OF+8JpQpnD0Mab7ol5ZzvJ4FDzSlJTWuQfRF1JoOHBuCvGcGBqWtw78Mq
CdVXeF4FS9wxwQgqHlXqQiuEUytFbsYrMIAtK6dE+wi6UrMHlFA2RmZaa3VswS6UF6vJCOLzmmKs
Xfvz4hkhIqzy0AR/f9TO/bsAyYyiMdJO65ABMREatJPLGXD97qEJkVqGDxQadu+9qLa0G4Uw/HBF
3OovrbAOl2EB7K2KF1F7IyRuG1kfZ5G4XvbWg4vOuKHs4OdOVUlEQSpfav/ob6ocopnZc/GDDG96
g8bGiSYZgq8Sieot9OX0dEhmGYiXiOkS7gSJedaOvumiRmnxCQ+snOtuS+N6kXKpzVNs0MROENdT
0BKijdUWKaSYJDu1drEpUmu6nDxOlGYhhto+fnPZ8XJjZo5xqQry9enxI0TBiHgFEuWs7va5Y5JM
0aQN0asQK3N8++57vec9ZwulNLOkt7UDwAk5yeomR36BokDJz0W+7HKuzhYGpBPWSOFCbPael586
UJpdKmviCUZQ2ImlvbtSOVdNH0+0ADm2xCTBBNN2Y+vstDrztlnt+ofJNhPIdrNjlxKlmRgAsm6K
kBtEby3NdxSclD9euHjRcqp+iPNtEaU3n5BAIbxIob9KIjIqR6/vC4EzXjfQq3OL4PXLVliHOKPn
nz9BRZ9uERk1Pzwcc6WxhKNZzJ4vOEu3aB59lWJ1wsS56/vK/97K3QfRICB4/IXko/irK2Sfo8RR
d44Z/MhcZrBR6rKDYflAfuAxh7xyKyaV0W/YdFxKfWahFzwv3I26UuxDgWqPvJQARnWT1wdySfCY
wcToFy+8133XQTk3TGJtUc7ZXhzp5P/RDFEVlx7Sq/ajX415PUL2Fcoe9zxGCJH/oRLu7AOWMk7Z
481pQUkrC+176zTU0kPkSC5Fv6/OK7a3pvvpPxbK5dVkKzykMmNJlHuicCsSj3ldcEyTWO5//OJs
6C+3Rx4l1SsRDD0sdaMdmS6XOSTDjWU5LiK4wCAQbCTC8qu29QV3Vh+OQMOAG+TzvSSXP0m9kfXv
VlWvPEqKUKZtmu6zY9CbCLQV5dP3y4Sn2SrWx2rfUvqdpZsNZDvcKNcvHr/dVGsC2798fFCy5sOE
y0acQy0be9L8jHDQ/jdjPK+qFmRpQGtXz+gxIwMPFETBrKxfJ7HCXz+wFvIT9lSMad6J1+wE9F/0
fhpskCqd2K6aSGRfwZjArk03PlF+gK7IPRDQhCPhZtGB0Rh4jJiaCntKud3SKVXtdQPRsFBlQZTH
Mq6f50Cd8zqlP3d/nbz2EX2UQZ8IN/EAyrbIp9cSWRNTcu2r+B3JtmKY64QKLXNlG45ppjXaGkQ5
AbNdKQGIPKFjMfXHzQoKB6s/+l/GXIz9SmYMeE0jt5iblC/7MrO2ecwJLYo+710dFPcsyKPgaPo/
8o3Z0OtNwg/VEI5APWFD5ZmOnUG2PE2yGV6W0R6aiC7SmbV90azBnBr3JrBl1Diaqjpvt8otensa
t0lo+O0+pJJ+HZwgMJoj1Adgcb5FbAUPirsKtHTfqm7+7dIMf1d/rrH+5lr4z3RkJmYPmYOkqbNl
ccsT/TO/FbjDcs8A0rBW+Ql796dgFQ5o7xLU8oYmXN1PTaIKVltfeIafGPStThRBQLK1ydi3tH1z
1tt5t4u0q8UlGEvA1iDbCMUr8rdXIsIlXGyBWamRT2tUVC5mN/5SZCicuKvUa1iPUYSpTN8V0daB
NHpDkewDhQhk/AJHMxy3sVWf173Vsy8DrTYdrCp8Vc2zLCO3kfpUAbPmN2qm/TWtPt8FF2MV6lMn
MKyqkqfSlcKMw+mj7+gUss0+i7YtIlrgGNzVCgJUsXkZV+Y8ZHx0mZYOvK0N/dCpHIssF5l+jUBd
yOD2cq2P4OKjB6hoLDBzwQAqRVY5TowRu2AEpHm+1KwnDei7jN6DeGxxlksmpvevkL3FuDNwmQVq
3t8ERPzk4vSv03Jg7XTWrfFBlII/DV0RItHAEveKnWZfGDOuxrl1UE+29VZ/cSUqiUDe6B6UACVN
9CjJJuauTif/eVTFQbcnI/zvfee/eVZ8YB+ZsQZ2KHbVbAK3l5fI5jOifOM/ACFOHk2vBAjWRRcx
/pN5B0bmpdGj2XUoYas8BmN+n5VYqAKgzyd3JVU5NlptpOf7HDx88gI0wo7xo+dYRbV8/bGuj49L
wG0fOD0c+PDj5e32neEbhxuaBAoSoXBqF2q1Na7MX+fHqHDIucRbXAbMxmPsxC/LDomF1wfMmmoC
LQp+5NyqzNICI82NOuTKO3rnqOTv4d8XFL60gcNo1gO1lvlgsu9naaSfQNPIqZpI4uhgJfxdqJMC
FUr93F3qznd9ZB12ELJqq8s0bZzhl1lNWh/NzM8aBKG3pcm9QtTHUQraKPq+ftNcpAXFc1PeIeBx
/xnjT5oD+yRA8djLUBu5F03HwnRDh6KKOzzkz9CqjyYPnTYU09Ode+vUvR1CXxkWTjJo3Zn99ybX
pxDZCP1CkRaJB2AUt3eikNA23FZWWusFoOYvbleMqFZm+0jURyjK4PjvKZxPP7xAM3E41wVcmlRb
o/xrCXA9gcxLCxJ0GKs/DiaGUEG3g7wzAEifCMKYfXzC4xkED7wkXWu4amipJYwbgwe8iE3Cneoz
e/05cdrh8q12BPNxVLcJ+DEM9O7Au4Lb+5xNPLBKNOoo4/swglJKJKLCcVm3NVic9abCBb3W9FPP
Jkz8nz9o8a6Bxx5IZeNqcrlg8j0X1skqCtftz8ZKKfkWCG2zWhWNjBz2xd9NZzH7pHoNkgUa/p9j
sOLbrebl8CQXcZw1N3LttkyYbgXyAC1YN8Ghb9XKSkHpnvnUp1dMGuzzKrqNcSbtIqqY5oT2kIDB
pYO5TQgj5iptj1St8A72O8ux4YAeCzBzdmRFOHmEbF59rCWAyzaATtSUR7OYelzBWMsnOp43jE/B
EeRtvKANeJ3QS2Fj9x5iC0IRlX2lFD9FK5ljZO9anBAqvIoCZljXUjM3NVFG79l7bUnU9s9RWH4c
P1I707+YiE1VYgEMNr11Ng4KhuXf99NLjIgsEdu35WoV6lHebZqLDDAmmTmsjPSDxuH45ZaGbHdB
I+fX4No0UZ/DQV8Io1oFldyfpEPIW/tYX6PZDkp2K04/zDTWeVLG41nw9lspTNo7yg5gE90lHEGV
7nCNkgGWXujglLAIuv1fdVs8HwQvSKVyUixjU9dBJZnnjU36gMa2RwnrOszlsxwu20giEzahnB9e
W1cTkDSNiFUM1JGavi4g7/iSqTdfDLIFd2lQl+50/MvgUJ6BB5cfcXYOYn8oLGklDmvum3UbGin3
f0M/HcYvwYzInfbJjnWCyShDu4LcygDIUEaCmrWsNmXApmQ0miB3+TIOeL7DPjjpPnYr98f8nuN4
SIYraCO4FU51H6hEGbjJWTkDYZljv5QpNqQVg9DogTWseTxcHwYrLxWtwRHb35j7QMhbDEUeqYVv
Gs+ViY8drmLCt7N1xq4DtzXcgVVyGeoHiwGx+dYO1iqzdP4vHbg7rNhekyiHctv6fLrNXagqDFOo
xDn4zodKr1e3adiTnp+MOTPfWom53MBTjUVzVyQ/7ANgpP10dNk02wMtNFEz+scBMSIftr3gPuYA
YdUeKGIpbqquyhBEBfdMC6QlzPPWChYDc9DUo1FXldYeRuZO8ROw/xYWrh2wdPPtfYdaLEZ8VQEs
6N3mNjJMAqHv+ddZFda5AtIEnAyW6yMuP5N9ocPdPWoLX/qZ5UHJqwO2azJB4rC8TOCE1pEJO0EB
XFgNBbuv/wGhx6KI5jznRUp7tQjmJL6oN/mOrQr52c1btpxYtCBLb1VjP4JJhcVbZr6EwA3cRf6I
qLhT8QSN5IQf2NkA5VjbeI9x9A6tuE4I989Z/020MxEyZVO8LoS5+1EJtGcQ6O31rc0XXodkZjhN
UCdEy0aN3nbuP6trcrcmnwt626jvrhqQslzj1+s+C7IvcIP+ecmIqOEx2H4Dj0eKd8YQ+s3ltKBV
02yRohVTCDpXQCxlnf55wOvJJUBOcbzATA12Szgve4SG6sAaeL4aY+EaIk3lITIkRji4uL1CLTNp
/v1bJzkgNxQZyGFrb6oChOBcoml+2DfOLrjA3uI7FLPhm7Bw95CcZbLj0OS/IUEKyRBrXGpO+o3h
67salADiBRQHCp3AY088j9nbyaIE7fUGfca3KJsv4ud9HnolaMCxcH/DBPYHkg4MOHkx1B8ep0Zz
tGJxaXP8HLUJQlnOgKrJZM9+QqrUjfbRfLxAjgb3gzWjAN9UAjKxc2SZDcp5I0ZxhkOlX1igX677
RINedIIv9/Lv0XaivvRt8o+m/ueT4Uw9O+DZZhRr2ZGQjwBBx2Dj3ocfeh9A8oPAw0u5K1P6kqWG
st4AkfpKQSAL9kfu346Ay6tmn/dmLN8GlOYaeyA4EaQ4m8NtJOSSborQ0FXPsO36SNobkH++553m
CHIzBCcOAZ0sTG5ibAAn5oMnvP7eGwVDCUszl2sQ+DXSq71nTJoMxepCi8kU9p7ResBvP79UmW9V
cmb6L78ZQi7vYvvZjtZlYMW48mFxdo2A1I5VKGFkyVkObpsghhDGeqZOO+0t7VvTPmcSieJ0VPQe
sH6Buc3EShUpgYqtUwMS6wWRq6XAP6mC1LAl0G31bMV9CIGxlDWpwX6JR+0NtKNGwtQ11rMfyqnq
iBumOaWKDyvdShDZKvxoz/sQrWXovkkEhN0S5+D+/p+REMzAew7fwahrTgGTZhk3l43C/LRS7RRm
iYo0/Ss+lo25vqrvhqSoNH4BCe4oYVX7AOeFJCvqkL6R/NMOZEsK1qw4GZYMCvMeyDr2SOInRUGt
giVy6+RzleNEYSyNMF/mKiOrkqjl6KNDRXL4bYufofwIitVbYskt487Qhj6mLuvCzbEMabH/DwnY
pNHMQjlOv3wRX6y2lrUaiPWMTlI9z8TjDERle6g/+Ws9A3CNyp2MkOux2n7FZxPPBzpsJHz8M+9j
qtQm0xRSsa+oURCAsthsGdAOOPiATvQqf42QKvzvrSdKOsWKi/9ELYX5InISJSxNrTZtti6Y1dKP
atfB6eocFPiDsuSIMqAd11MiQf1JkKUoOhGLj/9Ab3icVQCQvRuz59ze9zAcet8btCoKpACNgYMe
LlPyc5uodDUW5L5r9u5iL5GaRuDn5gWfgiVDkVeapVta1nV2uVmP0APLAVvcZmLDRXnSM8yuHXKH
1ezTKSX3HIysiD+sAzuVRY9Zi+zvZh4u29OvvpVHac/IO7rZesClaCD41VH+BBDro80ItGDWl0DD
00+FkOj9Syy5kwuK+5kB7xc5+nDnFDF4D6D+Nb3aswEJxqXafZIhmJE7hW++i/sZcynoCEX/mNSG
oNAstD05ae2EtFMwAaEnlj6fjvf9nlbYNZnPbafwgWXHIxz/dZ+XYNIeI9oWA8wiO01kcLEQ7xa4
+VqNOpGzDp8QFdiC31CWG44C5A2YSdSQ9d/PH7k3Tj/ip9FiZ4g86wJAYIGI6SfHoMEdPDzvp83o
qAHUDw9aZUqUAOdvmi7bzUh8fnh6Vb3cNXLSm8A8HNo/FCgD8P7UYYsXBHmHG5p1CB3kFzISUrlv
MD8YLCKhY9dzRKNXyIkIjRDiZC0AtKD6lG4jdlqP2qH79PmU4yJTEFOvwN9wFU0Y3nxb6CqnhaLD
JoMrd16tpCEXoWvjrkfovBq/cJo62mlXR+C2xmGHMOZcGFXWLGLAG5eCj715ez7jDEqa7n7259tD
xDVBhm+1JI6nPifD2KOGxAXzny/aqsHzXzfoijbQOkHZecaIEO4iusnGwMyjPnv/gNcm4DXgxxAC
woxdyBooV4oujCSsI+c90khXT8aPX1InYrq1h33xW1QS3tfYtTP58J0k6BOAJdEUPDzTamosP2px
qAzREr4aEM13yyttjJAqKlGpTE4EPlCeWE7BSt3CunXcu4KAtstw3zVowGOL4By/a2JJ/hvGRRIS
b6+5ZaT7nJzggD1U8gzz+kfj3q78SQlFOYDuvORBXYZ5D+DYy+3P1+d+7LHOpdySjC76PM18lTz7
JsRw6z9jYyMFdYAGf4vEQ0CSzV5zHs3yll1SSltH9RPrR7re19oAIi19V7uuzxegrBXCgnTMyXfC
9DbkwTvDFJhOweWJ9yNyKxyGe2q0bqD/1S+9CyTw9NpXqCZm0tyL1kPt2JDatlCyafR9LyGegP6I
oZbK4r/AkFv44cdJR4RSQJv4EfY+/Kkg1auAxxyPrNso4Ej/pjhsk813DSYkn3WSN7yqUALbSgK0
IJzYMJxsYH5UkNNqJDoluLtP2jS9I9m3UD02Ygf8+IixcAPI9yU6PtmPu9nwNBZ1ibVnk8r7clIe
F4YdXuYHsnotMfxEUDbK/LcVzSYJ3iV8OefP3OYgtLI82OLgUoqNrgPGLhey5xTzFoAcFaxood8i
tj5LPDZ+O/y6+Td6/kcI8NQYNWJQoDeiQmVuPCzgWO08UxO9CuBS6PjBTMdnkMfJ/zYC5vc1fobg
paKZORWe2meT4KomfEgKphTo2s9ps8UdhTcDK6aGw3kXzHUedk+F3vIgnclBxrnSfVcCZBy+/Eub
pQlUp8TFViU2x1nuxLiKwmzx9ByKVT9vuAVNtt7Fo99vebr4unYxjDXJ56WgTISk28ZFaUBDKr8h
57chyHJVMwD5atR/n+up4ccsrlUOtOlmtnXwjMF71t2oVXw4sLofoQrbaBViERFhMkJ8pyU2O8mZ
tLrzObGwCxr+FalJOAA9r3g392Sq7NzmyGFWCTHpsm2rb8VV3qxBHj6HyTa3WWARTcaGi/4+Ldda
n9Jdd4/HJfVrpusY8zqmUCg1iAEYqbIkkwoCz7AfVNi58xvRLXZ5MqJW3u2FxF/10VJ39x19UsDP
QF1RZCWQfrBYTMpelDFirYVyj5lnNq1zBcwgDKARt/0/Wxi2IUwziKHWS+qxzx506vC6+d9jRnVl
PQXDbJlKsuVhX8EY++Yxv7TE79O5uv+GUg6N/DPG5C63V8Wywj6Lhu4jJpAoTEVhSgwpTQK5qtgq
U5RzTtMDwLjU22fu0VMY0JaFYMugMjDwCItT0MG9MpfFzLzwYWzDupcKgK6twO9al8jcLZAp1xbQ
987AFOYFZWJFdzrS4Aqy8ZWDP5j9fQSLA6T/1bx1mLCT/fP9B+1L/8ddUyBergSUfIgnuA9FmUai
l6mWCLGEMS7Fk/uV3meoGEktTeFHsHOA3P/GLiEabBY7WLD6O62wq3nnfV+j8198aKscOybFce81
6BIqrsr9mc6z6+Pu4iB/QMdsT9Acx/wf/DtJIq4F/03k43oNZQ0E+ERNyynafesagBXcHEcJNr1l
sOWANpV49GmrkUEcYSWPkWCm02g6MvzMY1i8YeloRBMNaphGVvqnnxhXU/bDZeyOaHbSMwR46L0y
NDGM7UxNHyUNiHoY5IjAe0FyfzpZeVVDnWk9QHf9qkC0760mAK7H9BrDTSCh1j35XUtAItuNXpOp
uPdLKdfCYxa7YJleU+1UUMn66YF4DUdInvtJWK1mrY7/xQqtVpsGeH3rKFBvzc3Pp4KMgSTl8HPq
WVECEYLoaw1WqU4nkPhtqu3PqQ0gdfhjmZ4sJJlPAgapuDR8KgSvQs8oAkqgS7eloZs3Bvmk/u3V
t2MdMmK940vXyD/6/dkh3Pk2Hcb4qXbVNGRnR8o2vqrzVA8nd/vz0oWn/ujOKNkPhcmqxSFZAuEd
jWDBodfFcTIq+3XBK5MSxyd05Qedl/HdOurTceBpxV8mPeSZQ1db4aks46f97vcovhokverdnzmb
oFpDuXsmpwuCc6HjgItEV79/iFEqVP2WLo6WvvX4MQMhcshWesOkcicunvoxSMPcAU3u5ivwfEd/
IyRdLJCnouJQfl6x0R9z3QD+usD5rsv0Zby2/JuxVa5L2PleQw7T+rPoHXE6xrsitzQeevoM5815
2SceJpzQKycd7F4kiZZOHgdcOB40zvgBVY8bapIF41q2kTfVYN+LjQ2HIIySiFc4mkiJhRDHgkN8
HkMFIpHRtqHdWsxKmf5VeEjmb3chaZFpaseQvDZNtYTqgUST2kAQWoaa2rh0R0HE0d5iO5nB+Rx/
AL4pFLJFdheVRnXMuW12RIPv7aq2pK6Id3pfuFpk4fmunABPKTWVZv2hTmeoWvb9ovHfsWlrOK+S
C3zU9cbGCQn2gO6PnFDLAQdGntT7osFDpZjibajXcFfL433KfMOVtnghyPgfAaCzG6r3pw8hh9Ju
d572LxXYDwK8onaGQR2WmdVwYdjPTG1KcPRpI6MMj7SRoJf7KDRgAkBGzGd6dSPYfdiY8rzY46jd
HZZq6T0YqqCDuTRUCwHVm93DwqvvT1hV5Z0AulOiTOIKrWd50mBIQ8nrfSIhxdqYbtScrelk8h3I
U5lzAyVHI37IvcGl0j86Uv6MRKpBanI+/8hqwbRV9QrPR1k74Rd80KUmKeX1hMF8eFv6GcG0Yfpi
o+ycvYVn4mAc6Mt0PlNfNDlnhaonr8OtWWi5mI37Im7KF8ggc4m4YQXjhQSpStVUiMKyPXiSgrs/
WYRmo/PHBp24uMWfb51qzlTzM2Ts+isHo7bIxIGv8xj/zWz4iW/MUy3e5326dE5m7EQvhMLZMmGj
4ixUfIRBefMPsKuiy9A0UuJiml3PPqJgW7wI10rC/cIjIRKm8HVQ4mOYeQ7qLyDti3SzVwqwmXCE
jCFFzypedKnVJ3K3uW4bxqUGu6hLLHBBewnRJgpuauvzcPaeYKHUTUeqF4QhcT1DZbmn+6I+thdT
bLsC1ku/NXA/Bnu96fdhXEhkD6e4HTunKsrphBTIgZtjzcD96LOHoCaEO4E2KD/j2G6VJdhuq2U7
Tll05gbLbJPUX4O/n/r8Ogg2Ub8pp7e1GVC19hKFd0x12w78JQp71mEpK+9wcT/3deFkGzzuOemm
PvKI48NbJcJCEY0cVHmOPdzGKeFyelLvQbg4N5BAhh5nxLpgLoyunDEIScMuLVJUr7uNlPVBx94e
IZo4RvyQh72ehNJwzX2ViFfW0g1JWsnf3wwAh4v8nlgWb+HGduH2KJq8tNJR6FbGmqNSMvdCYXaj
YbTBHf4GX+hXnDSTmkBP+zXdqBYPs8e2pZ/1+9o8U0my5fm0LSLl4xH1oyFmk0WNjagVd7ODtTTJ
oyj+NqH+Y14o4zTuw35RSvu+tL1A0xGnQxx+fxmWgq9fyYjWAgwyghICsoqNdXof5yCvGqEtGm1E
9tOZt4KpymmOgT42sgC1/MfZmH4dcRKgHHQl7GZXRzinIYTtLlmpIBCMssD9H7rNl22MjOQwUUvk
R453PgWNY6DITICSLAuzx1u6IPnwozfNvJQouBiHnCF5ql1v5oIEqfxKa0UesIG/8WSNyYf6eSBg
kauMLGKh2E7NHO2KaCqQ6IqCpRyGSDX2zMvq0t9ej/aNdT8ND++ByH9hXKTDRC/H//bLzevn9p7G
tEibT5P+8cGKnNtP3EdtVji60wyg0OMgNlrP2JjsAyq/cFMUv8jKwevqGPqkpmHfKFqIFm0m+7yM
8iNRZ8ryruxwIHpx/uBV2BZ904PGcIkoK/sCy3XRWu3HRJgm5Rve8wxwR9J4I7nuSeefpXnxYakA
rMd6bZi+LUqIa4DutAKyYMd7OSQeDZpsqx2Sl3WFtMCKJFPmljW8hBn/+vn0vZoi5LqsGQDPBM7C
3VbVicZtucEtidPBD0nY6WKbveJnoeeJ9fHmI0L2dz5TGO9C0sCy2e3G7ZyOjXk7A39xGZfB1eTy
Vv2buw1UEeuzkKI1WzfSD5hRFbBPf/NuENTPF38tXZVfWAfR2TWnjW1yt4u8oPGk2xKwYnAXSy4a
/WNFI7eJGJ7ltfbpyOWDneINuSCECVGkP6tmx8xioIld05Y0D0HgWWjP/AweZt/CdHHUzbtXaIJ6
SzJY8+Fqsik3zhw3G9q3QP9QYRCGVBETnQ/PjI8BRkiTWB0hhpc0cG9cp1xHjqjxK5z0AafBPMbK
So0OH4IKlElL3We0bSHBtTxmEimA2R6kmoJwB6D8sQvQ/drPpR9r7Xrq36YE38oryGzMPhZIGLPX
rcCCneVggM8Vv+jNareddsr6DALw4yRaIyzM0vvJnPl01a8BEWpUZuzw/6rpzzfOOmYs/snjDtn9
40jyZIHOqu9nwb6hZW78YMqk2xDGbqOdjAdzQv5TAPp7YPcVTQSwQ3xEZUcnSlLEIJ9OJvsau4RH
dwPoxj1oW1B9Fn1sZwgyOTGySLzAOrpQWJwZHR8ZZpPoJ8biNm3nRTWBOAufnjL06T615iPEAsGw
3NX36olGtj/Yyn1wZd/MOuYALZhv4O0IafDbKyA6cL0TbWkLwii49kfq4W8K8dxS5rzwTETKQ44O
ovIjyOuHwubwmLufCISD9XJxLVwy6dsCA22NloZsEHVn/jFYCa8hsdqeArH9VXV1zAyDXM3RGZUM
fN8bNTTqjRD6NpIkuVa1jayyhVF3TqoepKIf+MEHE7ejD0JCWI89u6CxLqBoSvkZNib92e3c5Cy8
OYrvQhw0UVeKFFP/2qkqAvWjmOAOmZzMPfktGBC3eGfg5PIAJYCytxA4x+vourCgd6LuRMtdHLdU
3YNVk0fcQhb3AklJ+9iQyq2Ggm7Tg9ePxvO86rzGCt7LHGAFDCiI97Vu8KigFIII6ShcCvRcTRhK
w7WQ6lo4m0BX3SV0UoZq+p/Gmaq7ZU4TjTxVFBVRiHiYpeWUBPwmsfWdzB7h8ouj7dy+t07qyBrU
KS7VpVpdLEF/ThnKok/yKGe50Pgmj+rQ4WHWdKsrzJqNBGY3xuMU5NrpnKDuwe2H7Rp44DpcgSm5
4cjSiO8pnbYD9o84aZ/5eKvDekgtdAoJhQDNeHIPHsZoysIbeJ9mzTveQeGWQc6W71/nNaNalUkh
lxN4lwgH6jdsieySHi4cWdeDO7YPsGx1oWxOWUz5Ooc6jhj58SV36M4XRy4yMybLSwLLtaHjlySJ
uEuRVpy7R5TsArDeou46hwmTNL9J7Z2XN+JjnvBDCTJQc1n+Ew69bRzToKi3SkE37WPRq2HgR7XT
SkgESU0OtP15TaP1yY5nAAAIx5Mt8hIWTdOYj0GUJNQZIOb/30poXV21srSWm0LrpNGcNeK5ymET
8+6uMidICkIA/0lhHsp0R6MFAZV6PnRsBsinAEEt81OcfnjoERrjEC0U7VxwjKYcW1VGHoAGWpH0
wXKgmPOM+tQUvB+93rjdqhTUC5UR4StLywQ9Pp4Pmw4JmrZb4zdZyduJY9NZHHi93NeR2zlBWeuf
2w02eqJHFFUlfdE3AvBkV2m0ypdsBWjlf2Uo4xwLr6lsif5GsV/wOEYHkY4kO02cDHSYqY9BbKNi
ZFIqWtw+uSkdYZf2bxTLdDESAGHmd/Z8u9Q022e4N5nogV+P38EJvm055tDOl7wxvIgqQcc6yXGt
3aju/G4LcBWKQLM6nwPEJH2WgvgAwBWV9kNUaId2n67qwr5UCdxpgsPrSdfOQCb5dSCbPwtPGwy+
5Me8rTT6KxC/KBorzxapZkEy62V7X+PlaKAI78YuWiD2YJ9jK5gvk4DCXvvYeQjvoaSqbHa59Lj/
gslqsjZKM1Lf5x0rFxdMrlUwRsA98ufn8c2G/mqPkNEiQBsaIsIwOOvyRsJbU/v6FDp0d/kxuqxr
tmKyAfi2kQ4lj33fPJ8DsBOfZBBAk0DWK6xzYrFA0yzVHR/JlVnAvKRCod0yIiD7We1X3LajgT5Q
A+VzYQQu5GK5IVtYnj78Bm29j2J/JJLJzC+eXGBeeyUB4YsgUBVkHEu9BCupUyejcnCVTF8bDIO7
RnPG3hysjlHBiUR919C8kS8XP8oj11YneglXvTSTPW9ZBZ/MDFmrb4la9g7JWxpvyxITG/h7tXck
uh91mRWzOiWr6R/BBE9nz8Iv0WLgfmj80Ic5ez0Csw+lbR1ryX/jMdTLidIKQ5JoBY/L52+n5bfl
Y+KFslJ2urs1C6jkOJYN+rQuHOikVMapZB7hv1QSqtIhcyUsDLa6j9RYwfT6K14yj83it0XqNnJl
5PiLglfG0sZloGT1XTVwSP8ybiqP5BTus62/hnD3bWYGcUyHAtSr3GYucsDd6XhLLzB1zxP0SqpM
FB/enLh670L7iCpnEPgdEcbSgZJRibks59zMCMcqE9gF0YBCNmYiKtRiAFuc6fTOkW8h+hY6a00a
JEdaGipKizCN9Q+pHW2Vjnvfl0+YqvA/BMqkSnhkQ3Uz1B3zYAUdlN+ZI9q9saY6C67erZ7Y34Cn
+nidLcLyjyfErhKKIvXhPLMEmYOusODiuQRcwI7kTSOrrqYd2MI0za4Wrk+93WR94ol0SIwYO9W5
/3X5vWKBHuHtXDTzPCDmMZ38hkkJbQSl7ttDRretfVYEtWtb41LknKx+DZTSO/AcePdGfGIwYBTZ
CgKgrqOoGZcB9J9MIG/SvdvDZMu1TL3QgiXdhZjcDHtMOfAqyKc1bG/ctRm9Ms0j7oMtidIBcP9C
kTQBlqGb49goRy6JOflFd1cWP93ueBHP2McIcwgNC8Rjmch6iLKy4A4097lBZb5GYyaHbxeG7VMf
+WgR+1i7EtyJGlY8Su706fGMZaA46TwsWOX+Lsxi0spoDkXIxMJQhbWyddofX/yiQGkAIuvf50iw
jTWXr6gCf6EAJX7ZeqMViW2BVQKvrupnpBmKR7mdaL0lHU+q5wUlsn33U8eeIVdDCtukF2pAPUQM
ARmAJ6WY5LRpyOVOMHOSnVVPs5YV6MUV1y1zBNlp71cpSWd5R593nmOn0kr8cFwTZUy679SEdHGh
L7TSnEthmy/SnNLuY6/M0TFtLuFF3/B9KPW+TlDaiqs77HUfDPOt1G6Iac5v0J6zBH228bZ0rOxm
hErQrrsvU1TzU68RgfnC9iXYxYj8WFv+7RLiAw81z7OVqxgAHdL7wZB/n+RfZcE+bignycvdWooG
s6lr2AW7Rhrb5SzCseIb79t3KQ1cnQcWXQy1Vo0iPzllE8aLa+cTZLudqgJXLd9U+Ew4bevMuoD7
5aEqcmCAY+nct9M0S4fObTiTqvmN8jqAOXK90i+4stTr8ihNLOb5xy81uBAI8UZzrlH4sbtheSw8
28VfmDjyAWxfbfarv1R7eVpcIP5lHQqP8X5bvmhv6polxeN39mPkb2FEDGNQqUIgZr+IcPqBxFkc
1s/9megMgnY7ztMEN7KVhVMLr/KAQjDcc+7DSY7JxqCQNwJlKheosohx9iKnfweisNLZanMRiA+8
ouJLPWdY3Y33JJZaAtRqTNACZ1j7qW4FLOX+nqE8Wte2b9WQQXbRBwudNEKWdjCdO1qAq8+PH+wi
xRkUqlBJvPHJPHdc3NAtDWBUbDDfsn+8WErgxHZqB9wIHpd1GCzBRhIaZlAZg2lWj72CPoNdXH1B
l4/Tmu1eDqSuCe+KPU44B3MU4mFw6OKFmVvCZ0eAoXn+UZyR+03eK46z0nfaXg9ic2itY7Nzs5Ve
oWhxwvnbH6KvqakorvaJirO7FeU3+D/PpcdRlNNfgEjdJ4UCGmHoaMhWuf4goQ/O36hqVZb64USA
vALBLGfdNNlsCActLUBGg8uVYDiRjIDL9rHYzUcZWwEB6k2Dy1gZeFiEidNyYJ5jbrehbfskO/sM
QKM+dG6IHx7Et16j1hWpgRvgFAQHIDXzyHVvjWdAgCEZZLn2pLhKKNbIa4A62QE4aQu0FZCGqAxj
feCpHFKWH77gmpbG7euoY6jsPnJD2gcaLlxUw/cyfjoGSBUqhE2VTd2k7yj+lVM8HwZONS4E1+Vk
LCND+P6GiXnFX9x345F3Q7aWk09Qyyyc/HplP+lnnsvn4QD7C12A3CxCbKd1/k0OMqSy6p5EHAKC
yJogletv01va/73az0Gvhycq742UzTx8LoXKpXx+wwDpeC+WAQn4l7kPVsSD1FHL9N25Qq7Q0tkY
VI2gUu+TW0EhTPJbdeNVMLwHATIXrUv0827CeluzJJTTlz+oep4uup1r+nuVa2Cl5s9KAtCkvNUx
7qnl2mm6o4/XHRr97hGUhGpzdfhy+3CcZua2AmuMt/5TqdzD7lh71Lf8RCcBF/FaDrZO7zjh7bCD
i2wvMtNKIVjGXOdajecARlfEEKl/DMeG1y8UG1NmOP8t0kpPnksTFtiNhP2a4CaWrj4M8d6mQU/e
Ddh/X4E5kn7eZPpFeupIpW80uoq0cWGmqQt/d8ePQmw5dIQFsUJ4pa+SMIscwcFCnbH93VLs75+1
x3oHELFp7I3xq7/Nl5ZtHLmy0YKMz+qKWroNe8DscCQneUd3XQIcsh/Qi23xb1mBjoABk6rhfm4F
NKQd9cXqlj1LxzDUtPJPM73a9HmCIyLQYz/tC0s0Tk9w0CwbBrhqZRlwAY6qX0Vi58jGlWkbZfzK
4Sa9Yl0LHoaS41rUAChIZplKEd/9lyrKuGbFINh3Uc6jYzyNfUqH1O4ksJXK0DuSX/yA1wRsL2EM
Tk/lWWpSXpJVMPye+OX8LgpJ3p+U34eGdYRULCEi07Hntk2VaqCkaC7J98jYeYErg4zXaROkqZR8
1nB1y4cd+YJfqjb3G0g7fja8yD/YjhJDT9kcKxqHwsn93JeRZzRdH/x+++fQEHXw+MfgKLN9S3nD
nqfHmbSeoMdNS0GZAgpyAwx1UhuxyOzbkVm/nbAikRq98Qw+qx9n5iJSWSrzQP5e3d9eTgdGvIgM
OC2RZpMUlAQ9nJXNb7XuKeKj32kn3vml3za+xhIMHUCRJXy8OfOnkWzcgWhXlfh0BggEDmf0TXwK
N7rUYybdtQAEMypXGEzTGqJUYNXKou888MDkB//IXFLT1OWta35RdIv8SQcZa+vHexAOM2AVRIR4
NTXIJWHJiq/DdxCVtmusxK725VU0AT9fkYVYrg7qymbTL+EpQS2JUWsoC4FiFXzJV82YLHx5ulpB
/ATrYQATFDSyXYj1PH6idJ678wmYCXM/hGBV2vbMf3ca3XzWeQz8Q8JV2Y+lDmokJiZhA5wUz1lg
wB3JkSLW9HsynAwloxr7JIsiXAQJmlLbwh4wa01Nqzv0T/CCZEKKo5sId4vMowUP5h0I87aDyfq3
Efd4yMffZtGaC0bhlvT2V7tPchPSSUvHjwqZweFq37jDmo1Pw+U1JnbhseURj7FbtlDSSxa5Y6Dq
Im43fHd2O0jr0145JgaPsJ9sGCyOQ/kGqeNRCQWvVytd6oPNLEz3uABgRbePg/iTodknDzHVZenG
/macMKJjcZBXqMEDBvsa72T3ILvhG8qsKSOajq589wpiPT3Nr48qZdxm2NgrKky41MBJn2J/DJdr
ZsWytEpJmqtYBclRX2p/RutD8pXgiF0WRsFfcIIID1FTtJU3hm8/h5GONgVPzvmWKZN7U/3TPOzu
7Q8LX1kRwOxp5iF4bEf0WB7p2osJKgG9R8oqa8zfigweGQhszDFOHFT10FoAxb4Tes+nCSKfA1xT
nPqkqcTgEXAujIm48yvtvi1QZLIaCaR4txO8QzttkyaAKTcD5xSrjQLKNxJ+ko/ktCqHZuqOn8ct
ImBSVlUfLvR13nazqVg+Cm4YqkFNGjTy7plJYsZrGYNDQpg3rSLacUFtfzXKgp+fdVunXkL5VP+5
quU/+T4HYhRfMTdfGCH0DWnZ2f5DzZwjH8f/g5vT2pQtFf+4XHG008fjsi+deTnGn1/R0+K5Vrmg
xiAS/xsn3BUerJj/1LxWWJY17eh8z+o1xzefyFcRGmvxBE+iQuyp4YWO+FBZxp2v/n0+KZdKSYLp
rcsTx4d1uZKENPF9H9HL3uXukL8qLajiiS3SECXu5yEuHv7tyILRmaFyULRq7L5M+8L1cs5Mh5BJ
HuxQZYVkET7zodoyaVAqM5XTRw1B9BIrhprJcnJji9gFEzeos+/7EUTnBftTdmB2SHLKHeRA88LJ
O1hsVaua2MRlOmxBlgWWs7gm/RIl0qsshvVrz3xmN08iPQpqT1newa+UsMA+Q7FXj4PDrM/ZBXWn
ijpk6hthyHSaayrRZR7CTRkafylWyGePQ0FZmiApu93UvSmLKaqoO1pDf4dLjTz+pPCwiMj7b/Z8
ew+eOCBTo1QzhfmKVxvNF4YnYnmHyCLnXiRZUbiPH2l8oos3r5v+gcSdfgHgAnBArWL9HR7hHR0o
2lsh2DAz7CSppuSRadPvxTEukn7a0FaNlNXkus5QQYlKH9hhH6R2r1R6NIjsTtlvXusiNSlsqPON
kIN27BSm2Pi3wKtEX1WhNzeRO0jAsgVHZ/bkPT7OKCM57rEfmJ7a8ka8jk4038JtT6QurmGkCC8i
zkp1r4J7uFLHbkaohtylVZ/DJxAyQL/vhul4G/KYbOOhH3WCkNP/gSdpC15hn9cyhWKh3rVzg7Nb
PEbDwbp1WNoaxRbc+xzken/UrQ26EIIKPFKgOuR4psuAcv4+l1kPzJBsUhs8/a6dRVtdMB5mu6rF
+le3oeryhGVVCrHjzksm2VPk6fDV+ub20OqHzLwfGjnI8owa8t9vmXPWZMUoE3gosAj+fFby7KKX
HMRIjG5lMUgIbf7vnlPXemdDmg+qdLCENuDbK/UvusdA1Yh2k/e3lom1F6k9B2i5JTmyVzXPVIqM
c9erMNk6KnwoJbfxR8+wwTMvN+h6g/dhSmUh+5u2zcawMH3PYvBlzBSWWrQrxMylDXorP+Y3JW/w
Ee9wSESczyIKa0dUMk/65h83+9Kaet3EgBDDaH45pLDAa5IpU5kZlTEXW1zzQtqGNWEQN8HW/QkR
g9Sc3Zd9DKWZIc3JlLsD7ZX8v80qwpFSJCPA+THmcIVCFEMpaBzS7SqD3mxKYV78P1bECifhhM9M
3g0wHjQh12sjsrz41dnDPmzOzCphGdE5l0oQuoTVo/+jxyKMnLXi4bYEXUH0DEqMUMzACeQnW+Qg
InytQm4B855AI0+OBxbQFeRHij9cKZ3st5c7Y2wIq/IlnNXe4omt7eoMQKA+1fhVeP6Rc3YQv0Gr
oYmwVCpQ9w3FEbfInBmSv5KzhPIG06wIWGCLZIVlEeUINvEaG1c/1jcxbMfpz8m9ZKTVyfz6u6tA
K+J7QS8vjUbTr/QdGpCsWYxkMv4G/UPOiTttrEZH4kO4GG9QMohqnvXdZM1/rN0E9Pe6Q3EA4mSF
lInLLgV+HkHSWvP9a8vojTpDTq7bOlKcum03T6JHPVV3IJxsJKXClUqN/hqgxT+BHH4qpR2w54xy
Grrahne89uf3+BOKqph3rQlJUDBg116AHG1DgoQ7JPRASdaqg/+VdceQx/VIpXdiPP6OPpIrVVAa
uyUg8SoF3S7CiFWv6WQXy5QG5UDp2G5u6uNZvXyYr665nocAO3Hz2zX7/oc8fPTxjuqQpghc+qrN
T2RuAsUNVqajKH5UdB9nwkRUP1YjDCdc5qH2NGNKIKdypi3Q3w3+M3B+OuLFfdQPX9rTQR55lhjG
GY0EzlP6l8nHjYSAJawz7H52spTAhZxG7CwWS9MuIyrqeoO+Z43ooFNTJ9tMU9d0Y+1Kf/VC/enr
Eq3QLI7vDosU831xNq7nY+LbJorIzjIdegK5ZsNFsf3jOnL0TyRLqNtynP9y1K746eTZZ890ezsu
K2QP04qe496YxZq6QSCTaCxwvFmedsMXd8gMFFuCrdFn38hAYZdJUqCzuZcDHnuZlwzp+Zn83EEr
N1czz8v9+mq9now2bHOLkuQO5fAjiTmLpU9fFb/1bgUtczcpm+tG69RTP8VtHzTarMxtM4AwvYLl
C6SyZf6ltTtU+s6mj3q+aq6gjQDesuVJ5pYiFy3jDXLc5hsN6Q0/7AH9ti96UOMoGVdbWCnpeCri
rReQGG6sZhMFe+sxxuknbv3y1dV0dd1qDCuV0awGPc5aIW+f43E/NoZatm3keanWNPZXwV87y6VP
SAkTaXP1Peqqtqp6eEWbPsvA7ppam7C/1Ya6G0IINKKMcI/PmQmT6wGtLP8em49GztODU9U5O02f
NxwORU0uIWlSL5qtCSXthIyHeUBmMBp5NaCBD6gz6cucEHwnVZbnArUaU0QwkcW6iu37AbD1H2+I
CErLOkqu4PcpXG5LJRWulWFELGZjeOTqzkoajQYVQHyfcptLGDECXYXxw7TIRIpZWCV3Ki73yAzM
9gCCm+rhWRU7Kx9rvNKSJRIKGn5IdJ/9NEpdRFwA4VkHsTPPuBQfiIMHbo4SErcBofaKbHkGnQFx
Yb+p/O0+GCwDr47bnvglkf63i8P1mznOiW20YmVw5aQsp4QcUVcJKLZXM1bJixbwolCPkzlds8vA
4yLCB53ssLiZWw7HGlQ8s7+SJFRQAy/t0JpljKqADbZk8pkIRj6Wk57eCIvQuFNCBJ/S4dsh0Fmp
0UOmyh6e+zADUuGK1gbGarMIxCyBA80DaQk7fz9SUyKUsR1xmUJHYzw3Ce2OO/acbNEZWkZ5Go/+
lAb9gRdtiRX5vLvKnPt8iVsCY0Nv3q068DP2ARs0fAXOa6ysoiF8JRY42gL9KTnqUh3U9h0hvxgb
gUygKp31MfomveYGIB3d5yyNY4fcSBL3DYm1GzVVECjzm4tb5Ij1+ma+hOBgoHooo8MP8/2Z8aoB
g2mLs+J8YoXmxgNaUjlify9tFvB6mxe/DNSHkqElgXXiJo3Aj85ZqrqEUOmMsxuvQXrA0/hQy3d5
3RG/EFP9UDlq2IUqveUy6viCDbotK9Kt9iW7g9uRTOEUBhiH7MDUfTB9pSx+O/o2ZE3PHDP8tzVT
RdoSSMo1CjGBFOfpc4szIM4N2YAzCZpj+8Qy62JpyvmCAYhTXP/ZnIpU5mDR9Qgnalh+4JP7UjCx
wtEHTcSkelmAoi8zTgja9JYWEPXnm3tJh1kFbBg+JXW14xR4E8wkPDcuAgJkmJJrjInAwnruzXE1
wr2s9Czbqz5yjtNX4m5n/mmDO94uidJ8zP7DKGEFzFsXL/2jcZhGiHacLFL4Tn/YXQvFJBEpRe5R
eT9+a1Etam7j+6uU6rAaW21WjkMnlIK5mEtYwpMlFoCY3NlqVbUYczPAnKs00cMQ8xlW1u69e4XJ
tiGBSKiwOfkZ1dVFoes+ldbktb4KZcQjP+nFD7BlzVmXsTCLy5u0c35aR55WG6Z/wlRrjzBZdsTp
ZkYIjqPUl4q6dS8yo7n5CSYnFD8QyCrmAftqMi2A2m37ECqJHsoBy4o/Y9CEPCcex9UBw5h8UGE2
vO1KYg8lHfGpon/jUwItJyzwQQ+YarfhNoh9U6xzhuNpVuWcewvdTSRKq5BkgTQstVGtEM8WuCVZ
lUXscU0e0d3lclhxjBTiHsfDTa98A6JbMkhfnlnMOmpI+4ogmzG1iILWpVZ3a0wV2QVpzXzNWOSH
DDAnEW5Zcw/jDwyM5/GL7NLMGEJX3hWQmz5wVY0+kiQWr5saGcooW+tsiu5vTBvjpnJ7Ercao0UI
umDzo0MBWPvJxUAJ7cc4708o+RXRkVTtrPZ1z/Sj3FKlPIKycvKk/PE+LHNZQXs72dYjoY/nspIA
jnEmDLz4p7TyGCdmQ8U8mo0ao3+S3LIHdvd6rocUlDR/QLT4/oq9jffhRfIWTaMoPctUzckT+a1d
hCbbkFsZ42PecQZCP6pRqk5qIxXj0C6ixqDMWXzXHwhy/Ftz1BXCLUv9GD/IrLInQgz836HqIU+Y
ro9TaOByGoW8Z+694hRKMZE+5DSKQ6AKQQ+ZMUraPQB+PCO5svUd6MHpEKtQfZvoyOEnznYT2+Dx
Y/DCpTCDtCpTmFEaN53wncyDaq0WVHkA+xafxiq+pfUpgaNSxWb+b95JPRG06Fz5FEhqa2zSwgCd
tZ1XibdO3VRxUh14/ihfTXCPkcIFrKK/zxzAPWRyRz9LYsGu+q6VeabqJmI4rZJ91MmDfUIeNyG3
/adir2uZ+pAHYKw05MeWVWKXRNcucZ3/bQo+t++VRrxlklew8wKetgBZZMrGjbJ2eiwn//2f6SWP
Et1asQoMX6SI10JBaLbrW20njRUHDxrKDYSUqcGNE6OqASCVAzntf8eKYbVYIkLjQyWlSCRyya/D
k+NcYOHML4an1RUV3YSZF1/ceuktiecV+WKxrrvkME9rx9Hyun7xJS+VGUM9b7KQaVOiD+BZ1QZp
1W7J3v1HWHIZYFilSWLzJQ6c1Fj/PVaHyeAMy4DOPKeMlJpVrgUkQawWi+Fy1eSfuy7R8LVF7+rZ
qqQFETGyRftUSXWKqwgWRITxI9iv+l777TB7Q4bxcHGQ0iBXOEFex0GhzA5AMT54EB4Rk/bv9pHw
Y+ySw9zrkndpSkZl+HPVqKdUBZnpJw5ybVNam+w8F2JJcot2bFV04znoBkcqPxfyZDXPhhtykXnz
a/oCNPudwc45Dn8hxXh+tu5874itc4KYeRsLJnTkv3uZN+Um2Z+mzqxntkLzFXww76JM4QkMbVeI
Fy/83B7rfwzRe1Vdfpjs0wYd8QBlDgD7JbiUe3oPCkc6vumqKffQ0XII//J6G4dG8K17KjLhd5hW
+T5L92ziUUoGdYXnogrXfaGvnFniqZjRV+3J0rP2q4jVsBY1hq1aQIUkloPJHcpOJzXITwIRUxSu
Z1rXN0Sb4Y1Z3PvGt8jAPrW9yLFB9xbLHwsa8wyKE7iU1YuMXgXsSsgNYMnfPaMX3RgkklLnGoqf
2wvMptFlRrTV0Qr39VwasRzqfTQhLC1xYIC99RAuIVPeXQN4PFOOAaYQ7p/HzZuJA0WqQ+uccGzX
lfpE0tf6OTYdpqb0jdmqcScws71ovr7CUIV7sXCHLHdrLau3u34tA3nLeMd8jMW0ouvYhfDcpL5u
tXiDLBk7mr+lZZdQWu5oXEpCTHlDWyDg4WFCHi2SkdfewPremajC5eHrPkmbgBUCLXEqJkPr82bv
l9CF6zpqfXn3Z7N6n+30/PB65Zo4ieKqFs9DpBv3kjaxzxa8lp2mqwQlFFZDWDd+LvEFkLspYH4X
aIyJM8sO7CSijD9L9ylJKuDNszK7ECx/AkNYK9OZaWTHHGawQvsVqMV16OYE7TFFrOAMQu1FOxQE
P9i7SFMWz1/1/govTkMMSO19VHho1lovScF57CSAXM6XDqe+7D3n8pcw4Uqb945Lp5uYdsoHRZLk
IzfiZ5ta4bDmAN2OEFRYcvpuQU6BCxV9QeSiPEDv6Bamo/dGFEZ8dZPzFSouVme8NH6fQjCcw8fE
LHlM7pVG3yM+qckIwIWbTMok4F8lhdjsA30xOtw/onHiyfB7do1UMRRivT2dcNpKM1+tuUjXFBkf
r02PtEtKpR87/5QrolwIS4rUbJYEGQnARL0riO3nR8KH0Akfi2C9C286J21u26M7KPqWmlJ3FlO7
XBfZS8e9Zl67WwmTs6wNovqq8wQolTixDAq7SG8pvpqrUtf5/eJvq13cbZVvMEp4D6ETuLn4m6QW
zQwpFPDFoaJJgFGmQ95bg9L7aK+DpjSqGSc/zkZjD74TGc17kraZ9Xe9ins1pbZm9B34KG6jO0iO
holUXhVcmB5/aaRILnJrkxlf+JN2h2ooMCXRU6a2V3lmdDOSpyQ1YmXH5IL9w/o/5STyK2ajXs+B
NXvSglvpClEZhwZ8MP9y3+hS/4Qt77eHtAh6empnM8fP9rhHGLUH4muHHbR/Y3TvHa9E9JRpb4fD
wRTs+Kya08nXpHGnQa4dS+2HiRm2Klyunq0+nuwAFPVNm654Df5apZ9Ora4OO0Feb/SPCDbSCmBt
2/vNdTG5cautST+yBlsBU5a1OjOFjJltJr78y3rR7YiERqaCa9noZAv57yw8ESpylkHKyVpt+1U9
VFQnClQgJTitBfgf25q1rN6B9sfwbbOJ9PmzDNhWmPVUNBN7y7wiNSNLnZcibTb5EZ+IEgNzo84Z
Db0V+S2LizBBmjHpMdw9t/eZf3Kco/syPRH1jOE6QzTuJTGB/xeymjyK6bA/YB/gAAtiMQBSHEyP
ezUs2wG8WbmWC4IqT+/Na0u0gH0jPjPuPcY28RI83idI5GABHlKPn6us/fXCRJa9+8u8nAA3/ziI
6P2vQjC1Fy9LErI6pUU7t6yZ0B6unlsQH6FaldVSXbYftvXX2UEGzj9swGkDayyOP6akKv2qqdsu
3ikcJjRtuI/omh+hb59gia4o1XNdWD/vWKyfOzJBO4gMp91x0Nbni/tB8AreYJPl7TuMdvBXhpms
pW8I70JwrmPiLQNr6Pn3br7w0MPMnRlbm96659fGLZiF3RMtfgP9Jh6BadraiZUeT93kPaO9p4K8
TXUVEuT9ExGo6qj+33ApeBasg+Vru8Ar4LdiA1Hl/ib9opf5CdPK2Noj7a/18+dbIZ2tjMLo7cfn
2kk6xdggIU4IHNnwNoNcR6qLTGUjaTMRZWK84iYRWygIv3nilXy5gwHD+L6X3gX6ykDsrcGglSmf
BNMQdkU/JoOKPritvHxNw1rXOVnLcYIPN2YqfmgUgnbf37CbpussjyEPzQ32UvYhXRloGW1aQ5+b
4G/ReI1khZORHSGBM9G3bVQ97+ARmYqNGAQg5WUMsdBbHtL1y8io8j0/f2IWEUdMTuOZB29n4pJn
T2PCl5bSsHbzH8tDe5XCYsY0UnXEaEvaahLhn8TpzDYK+cr4xPDocQlbo0B1FUGwJxThZNzgNK9K
f8P0kJEe5XnlT8Oteow7ljbPH1i2b96OkYB6zaP2AeRTSuuUax2s2iuG03iDWQGEdfOCc91eKgTQ
pLMOdGNGO1dFtFNTePqd5Xc91imZbP0Eh0u793kimkfpg8E5omhFZujMF8m+AVuoALpsBsEmE2OK
VXXZs9mRE58Xj/D8tLzvOzDxT/1p6YRHYXP5i+8WL+Li8A1weDrMk8dgQHiAVjPrGeP87LutFEwt
/5DldZH1SXyMRMIN8utIHsDSX3BNoryqGET6HspJqufvDEU1k2G5JSxzWWMlsEyAlSMo7Q3ewG8L
3Q8B3x9Tnv940lhfCwTYjxQJA6NNp0mjPhMVbvaUA+pc3LpXnA/Erb5cxfTNc3Ru0McCGsYG0RWE
bRNNfthBdOjcNjGiXHQ/DdUnQtjDGFd15jyrfRaznLZnoX9C3xHoDpezw2Ba26vIZpkk1x3f6QHE
YbWRvM5Fb9W47gm90+6mswehqCtqQnnYSHkSKASrbzfCaxUzMeZOdJFgadPUq6WcoPJ2zTmZyA9k
R7Ri68gT6IjXbiDhsxCb16k/ynMC9Or4DyW1F9Bv3L0p48s7/Iqn8qy/hP31bZoAsqpMQ0Iu6JqR
zwKhcWr4jCiZVQNiQcVWPeuc66aUgzdABJZc6kPKnvt3pj1UrFnr/QyAZr6bcgUQMNMiQC9Uv5MI
yB4JdyCIv7V4qtr0vj4y0fvSj1iMCTfkE5mF20c8u+uWVFrFsKDyallfx01qg7fSVPtBz+ISiNUk
tBrhgJ9A27A6Hrl/rxIsFTVhN6v/EMk4hPnkmo6pxNoJKENHWevGKr+H+2Q6cSxfnj128wAybDbu
lO/PQ1nYw+JhmlAhZ4opI32asHd+ba3JqLCC/PbehGwXI7znREIrlTkRTmSf2LsDWcE9miGxtbln
whTohFfWVDa+vCKjG3BUixBfx8kNJOPH19gEENH0fSBna2N7V5yZNpPB91W/0ibPHMli7oQ/oMBP
LejlH5aWqGQk3/pSs/K/qERZzNgUSDllTj4c35pFqNGTfEg4nBELa3ikJToC6drpL79hJ09dTNjF
4vs/PsVmwB8Zsjh7iq23mReqqtJLOdAwK8APtXcbHGgPoIcnqRgwE2KGTXCQnbwtu4X2TD0jvQq8
XQ+aVcacJHIff9g/ZVnYO8ic4tvFAlO7tb+7woGmpBt9L2l/8CJuKl+qH89l3+25f9XW/DV8nuXO
OhPT0qCiiO4QLCAhsXt+E6UxB8bvrySqM/RQ+Dvqv6tFnOylKHnSYt+XwH74xNGC4fju4x9OJdMw
+B2ZRjfmZcwtshld7lzya6K+/OQwK9bmsJ4X47P4SbfhZOhrw3QugTm6zPsr6B563yCQ4OgC08TY
yJitd4QKWbl4W9//eEL7JvUTjZ1J8u1NY3ayupIBluRl3AjlgOPiX3pagaA30p1LOLfekBpAZU/L
An+K/3iD9dxxuOB0Brn2cWGZbrEEuVp/yRcykiFaNwv7MUHHOxQf8kc73dBSKRkQ1EIlaqJ7bwSo
DfUUgDWrgWn8fjYzUNwFPWqj8X2sOLZYB3mkSVArePPnf0LmVeUsn6JAUW+UG46scKyqmnUK9F5x
PmcrAfKtiwY2TeMNQsjQ3XTeMh5ilv0KtCKrnAXsNYBt+BlX/X3sEWdn9vRZKmKwtU+Pnx9cfYdY
bf6BH1aikYE7CNKAc2l1WGB+BE7BLlS4fycYeT1MoL6pKZCoNiyJx2RkmhW9mnF1IUilYQfiNtDL
kFGFgeFZUC1QzulsMaxYGe5QUrbkTLh2/axYJsa4wqAdgLWNdHmW9VRMzq+gbuhTcaHLBeov2WsN
muD+MX578/44rIGHweGve09HdYKoKY1CvcJfwl4dSavH7QtYQSKthrQwe00TbQa6K8m4VbM0EFgx
1LI8Yh0HCevT8ve9UAEqhIzAVW2M+p2v9o77MoszPPPChIxkaEGuti1FrIiTC7eU1N1dEbZsNlIR
Rd9jzjhXgCpIttXXoolsObweIy+PFMUcZJjW5qhob5A4bzTvNWteaUKGhof5xnFFwiIUbxTf26T4
vbQdApXG1K5m9dpAt6MUaWL7ofWwKYrWBnA30gd8V3PeDkbFCrCudafQZaheZm0CCzwmeTQskRY8
ef4vKVD2G2HMYC5UuISZlhi9AS67dMnC0a5tbL9qaknnd08sixXlyRQk9+Opb3hnqpgjX2WrdvlX
99oiJSVkBCzRP+4xnE3Gy3WOcLmIvLKsUt620yH9myNX5sehZrUvOW3OPs0uHwymy/IpBwCwpWKO
HUZSq9kucIId47ovEvEwg4EXYDRswJ5ncIFvG7+2qKgocd4fJlL7B2vKlsjJpjqDPr7f3mETHKWr
RB4i9oi/yEVN3fo9bgXXHYDbUAjjVeHLPoqnsPj5ixrI0gMJaprbJn+bz8sjcLbyzc9+CUc1aOJf
fhCCOGEo3qNgBpBpQLnwLmf/nyMiWsw010KFvfflfmJfApQ1r33x6K+dFqxVd9q4l8OEkj1AAkK5
JYFeFXGYEknKXkG0a4Dw+61WnmnQvxtSrgoVXcwkaodM5hRorjtGT2lyKFdkiyd7MVaUvoWvko0o
zd3gk1XFMCQBBoq3Okt+CpeTLYzfFUIFCG6a92sIBiDFtNvUO0Y73CWo9GKjFRRFdK0M/lglQNeh
BtIIhzTDh828gZWZwzOXK+nsGmNPGJtSAvx3CRjYn7zuctNr+6xJZpzkuYX3TeK+fOjrQjgncsrr
dOn5CfU/WwDqPzL7NZSEOlbh0k8PzTIx/GLlf9nV865fhnrMtRnY9/Vo5bm82tAoCRkCKDWiI+C8
wpR01le1/boHcLpIhC4dQxZVsHvOpTr5EXy8OVtcghr1dy3GJYhNFQ1fEmE3EExA0ageWLy1Bewt
qg6BRuFZuxPwChzGrJsK/RFW4QAJ6C+++cW7vvYB45YGjrz9kbe5eh6SQqzuwQtnkm7TkeTwVeKk
McVtZHGMrVKIDNNJGs20qQS6QfEls1RcfzH1jPJQ/YOubMnqeeRXx+Gk8hm4abN9D4BcQA6ZynMF
6X2qV3spI8GcbDOCd6k2CLSydaeaA8SgxTtbK/je0Oc5f/PbOmOY0Mm9DZVrNQfoC8kI4U4kXo9Y
MGbfxMKHL+/6N1X39CmQp2CcXARMN11tDxzq/k3C7vvaNbbUZmLbpQ2iiXkhPPXFM+Vz5a1N6OJm
odtvwdRJY8u+/nZRLfrk+W7rf+sSzXTo555afmVQUKLNU0+A3ifKSks1BGr+QCQX065hifLKxsH5
brGeGOzug2lOf6ZbZ2Rf1IvQjDevavWozjf51Art+kH8Pp0xw8CJLM/lNd8ZRUhJkTgiq6zhPBTz
T+OvHaIdmiRYjV/xtQaBcbCifM+Q9CaKEV0JvwlvQcUA+Kf/rr3dXl6Og6QWsfYxlC+tTBwo9QIJ
YSU3UTuA5peY6wuvfHY4z2U5YmUWhqdFy2wKohuxd3cQz2n0jYJUW5BNA/UjwsfuB6elQT4leEhl
NnAmuczaGR2Io9SYDvlamuX71RUeg3t65NyoU+mlGybZ3MlotW6BIn22afqawM3MI6g/zNNn2dUI
mkcDXn/089F0PLx8OUjNIJ67UH6UBCsmwXJL4NgxSg3KAROx+NKdO3vqS1Zyo/DiEE8n2P6gdx84
64o8sXkWXbKGkWsqyn6ODaks9JMeHuTRx3JywAJZZaNYIkPuYodsPcwIRYon6ZMG6aGfpnvse91x
RewVrpP4u3q926F1Sh2Xc+Md/yE4JfGo9h7P4tsW1MCVFDECah8h34DjJMD23YgE1kcsCE1tjt4B
SAHzXW1O+caPpbaqGCZeq3UOkwZ5q6E6rH1eNp3ZyFXvLG3YwmISLm6FGY7+hzGPVEzfEQcwKl/E
Ym9qVYm7Jvnr+ZLA+RSaOScvvnVeXWj5gIVpKGTksP9rljBGpRiz54jORVSmqWVGptdQIuIJQ2fM
YHI6obMbLJxQJOL/N2B5M7q8dNFHngpFdisshIXBaLRtHNJb2Xyu4Y58LXIABzuA5pirPZR5GAEf
2mdDFLmlYVbcSNrkx6zF2G5JEL5My5oZyr8KxMoq36KxBODKjpLTlUYdUEl/49DYQZ1Y/ba5BP8W
xeK8zqF6ZnL8/MmmCxF+qNZlxsGRmkfsMh+0tWr70BRdQios5/0oeY20qsRAsNeShpCYtzxl5+5c
olDMAg1+HWsaK446YWEKkt2//K0kvgIX9aYKIiFdN4tG4AsZPrFqjYzNmqP0GeiE2ddz455mv7OI
8zibZZVr49GsapyTpZnw1vL480G6XTlqQIFFutMxqck5XKT+iRjGVqeNtBdYfOCqyRkmy8HWlB6x
Qkyx1Xw+nSS2sRdmgBoSL2RoBKZdbKKHYULtvny/ScS/+kYby/eMNbvnH8B+Lc4a9bPljV5qbDEl
qy1dfdG4Ka4rQoeQHUAG5Ipr2pglyFHoK5j9CBCUTkkRzFl6IGr5t/yJfVNanbdXgJJ3ChAUPps1
o9/mYCRC86Uvx79xOLwMkFo+Ev5aKPnfo/XWIwHQW1N8NrNvNLy800nkwqPjkbyx3mhBDgWcqne4
kITQJ3uSZrdz0kbCHkSK8b755fxsYkOD3Ln4g4k+FWOVbDdzB/H4hOZ+LPIUhg3qTz29Xigii/Bd
Q5toJBPMPHSqElNfY9yhLQMinEAjlEMDRAeBd+xehCSagdfTcAHFQT8qhtHEikc7zh8GnifcVJOd
nnFBI2Ct3RWqCaZ/4QPukjSmS27hNIdbcvFQUHORhhqXCK1n2Kcbg/PhH4/JK79dgBvzB1gq0uvx
uu8lym5+YyKBoAXdu+KQwcrxznzpNDEBrVrNBw1POV2/jctaiwbOv84sjvFbdZ+baxQ7nxg5HwlU
RfZpX12WTYriBCMRF+Iv67h44WT4VOLeTeXdobUZ/JSp/gsTOBBVr8HJxrayk/rqqfNukhbPMON9
/MrxvP1FLHFpqcWfTtIRTBCqU3EKmkGFD2nSvYK0Go5CMWeVDwfdiyEmZUU9sRM2tT40r57fZVoU
cvqwfarEPOl69xIB9B51B/81lnUXbyaQEkWO5JBx3ZY0lz8BR5Yx439gRM4X+El6PlpD684yXJ44
3Ha3vNL1UoGeiV2GuKymfOIN6kAF+WwVthJz1nAxAGIWvauSOT11CleY3el4rlNFH7utWfG6uumx
JBCsRGHBo80swNm7TLbsleZTbrVfJ3tIpz3hJJ8G87ZlaDMYotxDBjyKHOXYQkUWUC1lVH+ALas7
0xBObncJjJq5cwjrWTNtP2xLqQvbC5lDBgY0nObdghSegfU4c1rL8M/ccquQ2BL21jVwDQjWQeLb
iZtGYdmTo/SShf/5g+prg63Nz1RzcyNhbji2YEZkgRVNMx5hxR9ZZVHodeBpQn6Fdc74PBaNzsJc
lgyFTChsGBYrtjworxfw4XAn1LAVhxSxNpoOoWk87t7JyBPElNuxPOVDunT+susQX8tws92WW8sv
Xfz0sBZzyNiv0k60carXlG2N1wJiBywPiKcxw+vfe6UotROIAcWTXdCzBVxJEAUQDQpEOIoLriLL
BebJWP0ZjqCAJsSu05bl4fHXAObbhcHYVtGSFW/upwbFlGwbXV7Wy9fTNrxFezxA8c8zf0kh9/+D
0XK8jswaqNd5HEGTAxCtVciLVExYkAu8gKB7ktNcPQOqJHeEiWuN6xhBSjgUP3k/vmjMfMa3J4+c
FOhLnXLK1R2hqU34KJWNisc5mzCEhdY8e6qjE05Tg0GAHSXV1tZVb2RzrYo8ccmkmNsl0vzPuf8z
YAjbwnTXPXji/W05mxyxpIpq+USP+wrk8CdmOTqejFaWjCQ40VnsFAwX/tJlME76+J35duwmxqq3
VvWAlkR5v38RzRh2aEI0NHUJ8lP47GBmrBp/TquRXFMZejzRMSym341EFiLk9SzhsFfKEtY9/eoK
UiYGAMu1YqDBFoCZsOjuul8RdjKTG+FLRwYmNkBupvuPzuj6nJUqWwUUtG9Oa6kdEzVlf0K4R6C5
CympYJFABQkemrjVKPLOA8Rwi+kPI/r2YKCWTs9hGpAgV2L4Ix6JMm28m640GnCzomWWWbnbZBn6
ctHXYi+lkgK153nOHiDFMEhkEmXpLr8kJqVXWFXWY059q/pxthqaf4jdaE4UZFw+LcVGGUqDBgi2
lkFj4fkQB7jbp8LsMY6Sdo0o8iQcIKeEEaf8kEgeLA7iSSpTEYifpouh2MwaCX5GubR0mSV/i37c
96vanh0A3AnC6RfAK21uXy45sRi/BRYEsdeOw/sBzlPOs3qfPID1rmiEvIW4F6Q7Tead/JSDn45p
lN1sC/5NzfyNtZ2+ZgmcMgXTDYkIZKxBXj3puhC8hc9srWx2EdjLrwr33lRorJYmyNaN4vbXIHe+
VZDBv/zD5T5u4n4raZke9t0xQ2WuZ/zLW7pIDiHk76Q2r1RgCPLW9+hvGiNqk51sQaOgkTjd1Np5
+nUFpUSJSl4c4EgqSec2dWZDZevzNuAGQHFikpN0UU6GsD6MwBNFbpexYbFDw5wmLYkcPTGzzj8i
xoyGeGi0k9AvJSGXm/3yzRt/i1KWj9W/L0epZ6SBNlg7ni/IjYYP+XFFjTodI0Xuz7Dv63cKvtw1
PV4PPVFfzl1FkIEqr6BrNlb4dbcOX68/g++DKip6zLIPJ3P0zHzgu872Y2Ui24XuYXTxqbE92mpr
yn6Q2/e4WkuJG96Em4r0XjueutvPZ0tViry9Xy2lX9mzoxu4ijC77ov9fJm1S7lRpbcNSxYA5pKi
/WkbY1+Tn/yFBiW/KdEHXb09M1EnUK4ib4ZtBB1B6N0jXMsXbqSuKW5mNWMQwVYuMy+i3UCWUyNi
guB5HgmHofbJhyGu+EQc9/wKWAsHKb3nOs5UdZFWfeiXh3PK6MejBflCpZVgyMq5wczl2AP9tNDs
mL41VMGva0E0/CzvbWcRBxLbxM3dqwJILOf/5H23pcAijglPh5Y9SYUUj1E4l3o9z8mwwCGlErNf
Hoq1mbIpwYYD0HK4R6SA5e/Is9GmadJzSD4zvG1NHPkaImkFfABdqcxY8pshTYfRdAuI4BOLng5f
cxq8o0DPCE7E01mLRn4ibIxHx6P6pTyfStrDGDvAE4MreO/o4mO4I+a3Wx6a7bqExASSoo3nROxZ
idSBprWALMb2iEkFaiGbRWfmR/C+dv2hyr66exJuexDfJa1CeTk01ueu3nH2lbF6LjXdJFxAmL55
ylaaI3Tj3xjbODoLVqv21RDO8b9sa2fgq0obenWBwTdVnxxI4QeoE8YZc8O3S1hBBIqzFnLkYWrK
MLM+DOB+nRZz2JiQoDsK2E4gyERjky0GQPi/R2yJpMIOUdYiwLZTInlvRXd6d79onf5wtbXQZffv
P2wSnWV0o50BLsvd8mTM2SBxVf4JYTdejkmRz6QMRNJfnwUVa1Ru0+mTakSmRYXItnKzxqItV5ZZ
6xs9XTYgrJgkwZzY5YcTd6LocZWOTAgA2ImY3TxTPdoCahIssz6pvf+KZHmTchZfAXrPLJ/pX3sU
1+g/eYza9TPcE/Bh/zpuf/iSR9BA/hBP/QKf7ZZca/gCWCKJ+vE0AYmfNgNOkPEr12BCuoTA7lvT
BczPMNwBZKTmWLbc2SFvMgYLqCuvWvGOgIpRC4/96KtULfn15bUE8TVcbIzfXjP3I1l9dUQhAGoT
gINr3CCBaGWWOeSHIzW25Y2I7095POTwuPc2wEPETSO8vTC5HfYV20sZwxV+EKz5Ck8PeTRvBap+
+lNXR0yw7KQtmAZ1do4axaDoa1o0lR/szLhad3w4aSP2Vr54v5XEZblBMUisyY71e+lIFz7zidmU
uOvNB31dd66feGA9ThBtrBhxXmpji9nCFn3njWdU3sKkPmDF5U0QE0V6zeb1bHaiTh12ZE1vxdhy
Oj58ehZoJjRdtSkG0N/oExfyJ5VD7rnQSoB+3ft/N20uQKSor8ArMSCWBvic57OqhGvusX3Md45Y
vhRZQpaJfVJVpSlTZcAxCbmAhN6USSY9WElBCP63pOYEDNokOYoIUEabksamyoKfx5teLakxXbtI
zfGBbRMqQpYpKnwWz0tVbDvqyfopuVgtSepHbiQxJxXTD8wK5iJsMOWHMhdISyTcVADFk5vnpgCk
JQzoRHVPC0RxvrGO7+zh+l38ztq6S5U8zDPDMsJto+sHRtleDM6nptfhYK/UcwDqFBwjkIxstlm0
Ihmk8Mhr5iQ4viYCafhQHwDUlHxrnuNTF35lZz8KiuRlPj6bvOyrWurSAGSscu1N+GKQHbEfKwna
IV3Kx4GTjVWJgljuTVJc3nUpHyu8D/1BmGDYXWhcjlbUM3CSjKV2mIhvwaiUR2w+0G3EZXv/Bcje
6it+pzS9K8CBey13gmbbicp7CI4GOuKWug9ItEUR2wGQCXwyMjyEFyInujPDxeoVzfSxsMOp1WgX
zqL+Og4H4ac1N23Hza9u0+to8Gc4mBhNz3Rpot5P6CnomRTdvv45jNfxqA/bEcfH/2XshL7hSvmk
SG6nI/cJd6GRFWN98VQsRyBNOyIsO4qnPwMAnzgQvZdy3cEHZXAYYIAfaGFSPisd3EnFCz/UJTQD
2B/n+ABUd5VI8wF+SXHJw4Qp5s6GqBOpizs5wgLEMwnRckJtu0WVyjR4gnDZtO2WOG7ebQYYHfeS
0/09Z0PNAIlT2miH60cK46jF29BbAWkQIViCi3ruRCJCEU7hvEjNtRl5wNr15wsPOfWQmdroJjEu
owkZ9PmNokwK6pMp9adiTah2rWVq4d2QRONdwHVdN1igcbUHjkVTf+yHLOoRUdkldBddEtruDRU1
jFH2+/a8UTDBAfddiKLwiJNbkedpYx2tnzDpmp+vdMBwG7Pfz+ncZcSlncdBRecjRVccS1GrgG5U
fywnbKr6s52wOSBQ3If11Jaay4lOXGDHPsPBVPo1AHNv2p2xq86TnDl4uYIPYqBIETGKzLW5lIm2
Dao3zfzRRLU0cFy0MDSrbEYT7vaN5/R3v60sdA9mHqWWHT9IB2B2Gl9g+ECw2/9wB5VPC37KB8lm
01zPLm3Hl376HDG3G6FejOZOWtm2KGccvPjFqfHq5MOya6c6CaChBA8rM7r3xcxxd1Ma8TbgKiZv
sGRmd6CQr85xzazeTQhypyMrjMNZ/eAoBiIXklE5Cl3Wgb/bv+2ubC3tDNf39vQFdivT8bECa7P7
SPRBeJZn2l+mnYjsJcA4AexknIFhBo/lJGSvoBf+UmjaIL4+1L8c2R62EYEvOXeNZnyJXZm1/yFO
MUuIn9GUCDsm2dwijYCoNfsopROBAr399J1I+KfZdtb/6QVZmV3zf3QfTDpJUsejLrLa2nV8LtPm
1QR4hDHl0JfH+J1Yzm9pM8UHH+ji8On8SSH6ItWo0E0T0qlO4a67HPSRb0WjWfCI5/3IHOlhJrLz
LLWWQzKdRziSdKOKcFkgqTtoL7Z6BbmZWfx8xn03uMzmqSlx3p4L2NxibdKe4HNlLggqKM/OVXkf
L/tcXsLzFVHKeQeppQRDLaUrb+7L/Kwyd3B79oxqzxlHniKzb3ZZwMkOBecgt4rce8yVR/KKd1DW
R2BIFQCYsd5bN5dlxdZpnxD9/aqmV4I3GUsmKyrjBSJe5wFdH7vyo0YS/kxPbxmCsyMBBQ6aEpOv
BNNzHCEozJ5bZgG81JfC4FtMkPkQVzdcnBxCnVl6XGtgTlUaN02fcoqiy36w4gZUbTzHEKsZH80N
lLUURa5YoDKDbyRYFDweb3z/HJDcbmzXIUs4inLB1UB+TCRm5jz7AL4n/ma1Zl6bJ5uJRrqkwoRR
I+WgtyEAVQlZJ4R1jHbDLxgTE+h2q9RKrNgCZxIRwyEjNf+MqNMrhEEoFpTLBB9FiG23VyOwa+/c
MnTy149FGRk53dFD+atFLBCWStiqbIv/S+eMe9Jer6pNN3DGl6Ck0EtLx+Zl1HiTIEZ9uli/Dp3O
rTNY1aadX+kVGt0opg8oOzlwinabSv7tycrEX+H2DlWuTj6eiuRYhHfxSTmroJguEm5DVq3lPm7T
43a/Fh46Odbu0J8m+swFB6bqtTaFeM/z1KfMVQ3gVClimdvAEunaIsWl4ZG2ipVCIxCIRfrn7xxM
+ITU0XKpH2GkC6R6alThk492/1epEzRwQi9YA+xLzEbz2HlgoOzMd1T5PaHF0F9+Pac8AZ/lEW0t
5Bsquf+DMNx6Y8uBEfV4FYhjnMLSrOJD6vW5KH3G6cmQMdWI2NMlGyJiSjt2XfRub092CsQMAQAv
uBanfIAKqpgsAPHrHh+569dmrvapGUTFhFz4C1VMh1j0WrBTDmmFb40s1zsPWxm0XtkoTOANPtyc
y8Xzi6R6TNvf29QNbj/yvtOFQFMnzlZ3w1uKfr+S6dZytzrc2H5M9Tx4ZZfqIsfAQW1mETNbx/mb
9wTyavNSbFmfPWaeqeH+0SUzzOien2K/rUn23q0qI5XgQXOJj0pzAYumFYT+MRknE8YF68jUFlTZ
pHWwn/nzUWcq1IxbEJyTPUtXJnEIcgcvsOT7DZ7o+nV7UKovD4JdOUo69eqJ5GhNU/HyZHRjetfU
8xKgcjsMbDEiUzTic+R4G1NWb3NvZXaJ5+hQTisd9r4IfBTkTBBGy3PDECjzxEEnqBZaYZ/PdiTa
my5VsrvTC3I2D91lHAqbJuf5lJXEFF+vDts4v2IzHFVNf6ugwYkZRQr3WJrDQYxkPFKeiaKy80Qg
Sn9FNVUTc6XkoxuYPSno1xHtmMn/x7o6jlrZ2TUR91ZjzrQevrwQ9iBsI8WOFVE8jjaeIl2QyoTv
neYtg4QKzu3K0DRSAVlp1sdcd2r2wL+OPCiVAKU+EHjqjzV89TBgegrqcElSm7xFFUxJVF/KQHIL
P+ALBjUuwpl3Qtx5azAt3lfQo/5o1+0BeoqCUCplm3AY4g8DbMvMAaGLViC5slTMniyfXoYBb+fF
1xThR86roJ3zKx/GjFe5LJcYX/U5gH7D9axluY7JS8ZJcIWKmqOsfVzngX1TOaur4FQ4YUrgYhWi
T/KyEZ5/EoPqZtTPy3eoGgUs9YNj1Uo9fA1AuliOufkDfIQaoMYDG7aXEQRIG53G5nCDDq17fS+B
LEz5dOmDO+6CIka4TJn4ModlZcffY9zCXFbT8m+BN9wFScS3Zy/oMuijHNCGF4iE8Y+EVka6eKaX
Ra53M5sXXmTmW4+o2NGvh45KPnS9IqsAMg7epOGNcnn6zz/ZYKMVKPtnvdPGX0b2qFjfWShv2gnS
AVZ6JuFbCmPTT6QUuRFvPCVEz6l1D57XCscE3BDw0P+MO1Ol1JR5l29E0ASSuVyiidII5oaoTtbh
sjszslfAdIyvbtvKyjUO2Vz8coavLTnpCMgkbeCM4O9cAEolq32WEDSE1EDbV8CdZY6qfLW4jTLy
LPtmoXBM8ofPov4TnGdcHu9KpA5q29rxTrDIZn6EW/DLYn4ZRa4UPkrBisJhwV8lENGfWJXMW5KF
gwMW1g8EgjSmn1uMhoZyOveqFG7kZ5g4JNdmqL1mep7CbyR9qUMwYauTNledQ3aDa4qzQzI347qn
e0j/JiKfiT3/6MXMD3YNpYV3t1AyXdkOKoEGzbMh6N5/nox5FfMfR6xjFTK9yQJaomS5p0Pt5Tr9
EkJ0z7G7au4Jb8ikCuW9iEnuzs/Fji9mrhUaVvijmxD2iP9zUAOjwaKrdsIJfjtCGzG9WSiwgADY
wHOuyL95I/rBAEhrA7muwzZHxeslvZVOwEFerNsJF9Kem3RKf6TSFgimI24ZvfGBZwS6QFC31Mzr
15tbzpk4BI2tPxL6iwvql+ViOsXtKJ7XtIqncPxR2LrjU9OlzDwF7fei1fY1hZrfp+iMAbJz37Ob
PQFQs/Co2vCZWave55115GaCdO1jGqGiLiagMGK/95thwYNX6gMmlKtv8Lgj6TgrmQHGX+5TMXwW
ymPSug9UyT98lFe+XOKiFJctp2M+N7bPwCnUFqu7lejbNzdtYJiPPqkVrXKEiRzIMJ3cX4xO0idW
bVpR8fnLZOet7ILpzezrlsEEs+vNfnmjN5yGPUD5RLGF8Ccn2kJquNCyv4+pQ+CqaysN9OgEhg/e
X1/8sd0/loex50NfzKSAWrmyrKlGxZu3YE6ugS09H+6IKMkNEZ+287QFuRm2SsXxQ50S5aauveaz
7vJzueZtY/d86Xeor4zwlxNqp7B1FGlXXX3eoEwXGwHcXDvtyai1ImtmANypdQ8A/YqcHjtgeZrQ
9uOjMOf7Jj7/1bxdxQumA4Dw3xjAMFpvgDqZawjJVZqXk2sGm5o4jc3jf4jSlHEMdoCE6EGAsHNj
UsRVdw/rUbW0ylcCfcluemUuQGNQHgXxa/HqeWm6DiWzLMsGQhUs4h7CZhm1Q2tA6pRkTBTQENxa
9F+QO+dW773wPxEoXb3PtTMgijavmYaC5GRIv4uqUJenQg2j1F1w7pXZH4jM0ZV2mmCo4vvb4uSV
lbJQXFJuxnLQNJvlo4TyZjJsaPg8bpelk4A90l7A3lowsx/YtNiR5x10YXQizh1mmj3e5TW7SQ52
DcXn5zr45GJ0yto3XaheZNWjQNbnOFcz8PD9u7QazoD8tl0dAwaCiI01WRuCClF+k3o2EkBKagoT
6Nj5utG4m7PmWz9dHkzwyRsbOhnIEH8LKW5zgiLATVZZJA7XWJAJIxBT+k7S2vMJzDjIp1HOS/q2
r4Kw0KJHcMXeX9yh4i4+UCwM8xdde1Sy5Il7k0e3B0G61tMmX8TIT6kuWxtzvzRB5alzq+HbOxcw
7NqlOYsRsdyg86hXuiPuHI6fUzgD8Wq1P2C/ZLlFtq1sXmW75V+wU4GjKA+9mL1p0XUVAoAwrkp4
H8OjAl0ilqI2+xySiw81I184BLX8o9hFYz/gNfPwrUlVF4rtP1zbMbb2j77APSIlEybyh17fqXcu
l0cs9LWgRwBWq5NO6xe4TCHbzONbAE9q55XBIAP690a2UxQoe85wBj0TQu+d0UnuM0B+1afh8Grj
+JP2DROTuKmFBeJZ6op4TR0tJmwTxGm7pCN5mHFKixHgtQLeN1MAdU0tiMgm6HrHrCLvAWaswRSE
17EheAhSUQwAEgi20bhuV9cQru5UuPzpvMJCbn3Vyu81Jevvat7UAfA1F8VDrar8Qb8IZ7Zwzh/Y
TdBS+/UAPkkc6a9qc+aRvkBx0lGAexNLvJBxwb5laokBPbBYd+NK9acSBBM80LQu6a9xQ9dx1C/5
8OovKjDsxDPI6MmhVUTm83g6U8ludm7ZliQR6qdAPsmfWSjUOHsX55glCgX/fnGvecbiBf7a1odS
3PCYjtVZW8DSOJV+p0r90lbkvpgUTbcT45oRqE0EAR67p/ZYfNxmWQGV/pNzF2D1KUAGRTGX+Ttf
Up1yMP9GEU9J4qr+j/ICuagNKHbOlnu67LRxvXtoofQS8R9JPFHuEGgY2LzEnYOGmFvSMdm6gqUF
pGPkYSKdDyFBv0shTDK4U4fHjkk8pcyUPDQaRzd70TNAfflehqE9XQchOK244flGOksPymqNttKl
Rgoi4WBNatRG9GPYCWQ2J5uTPG0796ym42si/TeWrK7YKMZ3PtsaqNrHkCekQyr0f9rqtxgbyitv
G1o0XR3iOc6UhVWRibM+J5kIWARp1qyVRwo31wZKca51zvpdJ4hV2v6SIsFAAqxfy/OAT2S7SRNZ
BSFFvxFXgTy3UpuF/dnpV0RAWttvFGO/6ViFXoHB3PaSX7kHj3U52fkph5B/FWuZ84UOruaTCasd
hd1b02clREis1DgLaX2lrKJNagwfY0cUbz8wTs2gAjwnzZolRASiCf2g+VDn4ULfndZffJBmmB9B
Tyf2EaV5X2gxqB4v1pJAEOUOchIPJLIk2mNmsKA8jMrZDpJyV2dWxsZ5M2TWoaXClw9PPzaYQXoM
iABKcNvMolbZ4a+CrGIMYD4t4lVoK7OeX2UNHL96Mtu8lPMOOM2EXM+qEEHOvJtKoH2mIygMiNlu
YrI234XdxEDmwmOzAq9WWib4234dQktFr9hk6AnWfJ4UYgTOF/DxsRXXOhQTYYOtlzvXRfu8uzNA
t1LKZK/dVtzhXk+YvG1TDHv1ZaBgRa0Mrfe07Q5hKrZISToDH4VJb3EmOGI4hFAEM0PFqiCx4WOs
NbE6+btgGmITN8ffW4TjEuDlJPbk2aDKLEqMLfm9OTogHjRNm9BB2z6C8dvrYJluV5WozGyiTCu4
iyeMm0TLkRjt8yME1r1XP5zVq4sp9i4cHwGMcAS/abpFu87zgM/rjap9PaO59/TaPUDYaKKTETgA
VEyLEnzm1MvOrE23SXULe2YC2prw3LuwZ80LcFWeP3gj4j95wUkblAC9Sb0+o9OR2GoD0BLVZdTs
FvZ49fNRzaQ5YzrMBCO+NTR7vOtrLYUC2NPWEntpTapnjQLB4MIbilDAmmvBw7w32U9h/dmTXdfN
NVM7Iwm8vm7FQsZBq24Z5HydbX6ZFkvr0fHW7n1Mtb8dW/X3gXz0TPbuyrrlSlSsJtspVBnEORi0
UHBXekz7VIWNlyjsexf262ojYRB47z01JTq4o1Df8BPJu5a+LBWzgwzYvlsKIejl6NsQpAxt338C
b7SiYo6SQxKQrx4tIL1hlsMxI/h0dj2pJoJSuo4xf4IhTiXvR/YvUiV7c9Z2HX22MVSkGDplCCwt
I/61iJW7eeJs+kBWDZliCX7KnjrQRXXLK4yTk1++Dvq9hkFziD5DLljqSJSWeMLDMmd0uatvlQbQ
2MyL+ZTDs7uDnZRkufU1FzGKXhHETnewjGG0f8Rh9V+b+/Y2cHyUQZh+xDLR/KQg5EJx7sIp06o1
QMgTvWs0Cw5E7K/AshCAjjITHNFvEM2fRd5++59Ir3idwvIl/6icInbt6H77smezP9thrDIez/cG
wCvHW/9P1EHGifaid39Oc3Y3MURKhNP/H05aOJwU/MUzVxvyn6rhL63mEXqkAWpPj6VEW7GOD7kS
xqNFepVVl6I1IKGVbvKLtAtpbgPaAt1m+H3C1oSquk9iXmGxZKc13VunTkKOa2z0Lt5SmCm6xbJ+
EDQisLhoG29YuU8U+NqS2h//sclo54f0eYWvqCixnL1yJlad+Xw5YMzBpUtRE0cbtdFheyAyOGmg
40uHqzFpGRgb9X0xk+mvQuZjcYemPfTjty4xYh7+7fHwmKhpnNCR9V/2GLCyi4+o6CRPh3Yv6Z2S
6N/7k9uo4N04LkCWCo/m7ZFwIRE3HY8y7A9WrCfhXavuErMiS+WtL2l/DsAELKSmi852YmeDv+Zj
fRtacBH54TTTpnGzRcxv7AvZnBnBnedEjsQLVbMGTN4h+rsyxmjjBMX6bqUeS2symR6lr7YOCd70
0cZ+YJNwDm2TRlakceOZ1RlCgt7RYAcvFvpBW39BVWpwYuZmM4X+Pdr5uGx1X9cdD/Rt4dOuS37M
fjxypwcalpI1WRVpcKH2dmOmoJ0NQjA7JNJnkMRJ83xmxfQSVBD5bIlyZxYHlDyVYzm9xOob99/y
eYHACAu+QSrsb709MkYpVXonWkjFagqXXKZ6uJMHQBIxhfE9+ILQi2ZU91rwCli/La0Zay82lmhV
NByLPu1t1HlQz+terPnKrtJBQME2swy1lSRxV3x4bz5Do8TnxvFH1ed5G98TD5niJEcJft7TGXfs
6QLjMAr54zjHE9TELOrIuLlMGGg/zJ4jwoBk0tiRY8jvucj4/os+WBAmZIsR6crd6L+4fxefAeij
zoBoMaRCNARx/x5xZYDr/YHJUHrXTKUZFzj+O5PhBbWz0RNnmV7mpAHh3OTEE0WQ+EhsqxGR/SQr
lD31tWnYSmxC4l9/21uVlFMsW6wEyOc9yF3KhMozOWtXqqr95Cv0x9VJqAR5dmPQKgBcKpIxSkjG
FPy65KhblWY5LK7PTh0lHAuJgcK1rX4uBAuz2duxN3/uZXVgove5Zm33y3dNT9u/HKxEbOV6XrsA
Ag6/FATpsO3K1ss4vSk3rFAui9jtFxCywlgtHDgE8Qf01HKBOFbqGViGurVgRx6zprfTp56I/AxF
y9XFDOwiAebvi+GK/w54yv/cakRCuOU2kealwt5rQUhvAJ+36pbXE8KqMB9S8sQzSEmOWcC6qjqP
sbn24lOot6pM0+n8FU7yQdQlrY5clBbSrI4ODht1tmI8CHRPBRj/yIW82KFtSX4M9Z5b+HYsXJYk
NmyW3rMPNfMUI2kCFAMmqmeVynSf4/Sk4PbojYg3ZIJ36csZNSeXrw2EKUyTK1VDoCNIu7XN5rFc
cwFsioQIFbvenfgcN7KxIT8bda9Eap7YNMe2dtTh4/n5H+LKG3OsjNNU14jwYxcDvxOIQa3xavaM
bJ78l68kXbItjhW6hjjcg/x89TfX9xK8i5g/hiWYikBWsY73t6X/D503Xk4CEKsBzwhlQbdm1bwL
TCr2wioJHv4kTWez1F+8rCZvVGs+EqJLR8R0s7oMqUzTwqVl/iwF09IW9povmUFkD6AE2QHxNeH3
0srEy5O3ecyfm3K/odD5HFmBNuN7au+yFdd/rA+Q9ul5T+q3cgjl5MfbTa/wzhAnCzLYoH7L5o75
fSwpTiUGT9uoU91P1uIm47oEvrByjZoGTbijzqRTWtSzWnrxMAmtEyb1kHuRsyQCfX7k2u609cYG
3K//7yRd3I2e5CWjTpToAUxHNS5h1+hj00DQNobCW+4jRaFDVcn9UOE/0mshpn+OCw31qzJd0Twa
r544Aa6xhVB4Z0+uXdPl/H7La28E6tx2ozt/ioY0iZWaTX2NE26L55FMv8KEupN4na09HaGewYjw
rL/GRTujOTya9m11hI8f4QUlNBFF//t9glCqK+HT4P26iYgoDPsS3ih0NlprFWBmKWW0yBg7FP7L
eMGmzQwhfpfufgsXjsirWLTAoL5yiARRhrsbaP1/Od2Uc6w9lo8qDLeflCNykMoy5miBdvpKiU8i
2JgHFtyHt3le3Lkdm/MQO3q6DSxeqtA0JX5WyP2erITzadkbNyUzWC9mROqciZKEyTK6+sd8y3K+
IVDGt9BinuCXSRj5oS2HZ9bz+bLD7RxZ4ZjZz3Cb6N9vvvAOI3OR8yftQsXfVpO884KLCUSGAGu+
p8InW6arF4Q+dCd0A0YOM57FB4dXdNhEjOQzNpsJlWGfcW3yGSBkx5f/eVHW49YkjZrIq5X2O2l7
L+A47UECnkBjcNBhPN7HTVGR908ZXBvVkdIrUUOSBp+99S3gwsc4cxD4cuSfQFJZtgIjNPi7kp9R
tZKcXAaroEEdNXmIHlF8WRnAqNafQlrDhyT6AgE781iHaLAoexUsOPLcIunhqFipMqo3uyL5zWTG
DDBfceq8fjF4pYihRtt3LBLlVd1YxnV/eMrZ9kx+RtUttNxcW/E1qJu57EYJgWCGLINyGdifr38z
ZOXnM0BaTRUWStgtn3QKDr4YjJ22MrqvnzFAwahiuo8qdcD/6exkactK+EwvHVVZkxiJ++UIMGKk
9yNC8jfnG6yzF+w38+p9dZd5bNgYXRuQViEFpHyTrB55BWSF7g3DYbyY7TCHWTT314ksxO7vKnJS
0Z7mbR15x8gEFftEbHjSAaTB9hs/YWAXbUXAYvYaNL916rwdGDYz2AlUnSJ8Q8I2Q1MrhyWiioG1
l0kb1ziEqrGrBoN1qp/MtQ8Dr70jHL7mZymsgcgLTpgUrEIhT2mLGw4h2NJCGW643eBtdzOgc3JO
FzYnC+tjtj6K2cmO6gPBIZeO7CWjWY8WbfPk1iq8NtraZ8oJxIXcwmyhEpC+dEtp2b4vYnP5EsHj
RZpkOyaYmdyT6HubF6xbFGWsFkf7J0yND/1ecsvZHINJVVrccFiuhBYa9ljbUyZLuT3QwaJjsqTe
Gaq4M0uSC7DY+0fxb+jOz3lM2Mc599nJDoa8yq5F6+zZhmfXQGei7mDv/V82CKFggYbFpnH69EMR
T8ADMdstbdgtnvZreLdMfpHRxDPJIimouBZdXjmpZmlOfk7aMDpbcmVT6LXsznZq7aVJhSPmITvx
bX4+zlyL0g0104YAGzu3+LXWqtVABYPXmYmecguyzwsHIqF83cJP4qvj7St8pZwcmXM2g3sywYWj
BwV1fwvNoIoTnM+n5ESlBKvQxAc08RfuVZ6QtLUnQ495GloYlU89zfPX1KSLqqdwQDyXTMO5z2y3
NBuvDUDmD/Lz0Y6OPoIHkV3a+5xGy2Fh4eYWEEKUuAlqQ+yN+piAot1wt2flSJIB/2qJJso2Fzkb
Lr8XdZSjsHacJK0UrRpXKy4IejoMziPf8f7O02/DaRHqo7jpUM8qNycvP9lWMcDANuInqCaZqQ5o
Y6iBnCpYT+8Z8DLQZwoqW0xAzgrtV52QC2ALkv31A/iF+wAutORS2VKANyUrKqme3lAVHKGukRSq
iGReJMtXRcSrKBxPHQSPCQAPLphOXHjcvxAY4hRVpE1Npn0TWL66tYgysLI6W78O0pj7aW0IdZf1
ZeSND4gj2jqd0E5uje9tsJ/c/jwAUHukdIGx9/ZpjdDWGafi0k7ModTJy6pfocy/YC/NDzWMP25r
mulJe73HS7dk6+Uif4We5XMCupGzk/osuG19Mmdz44JlHCSp9NBQJsSd9SrbTemsnTGWMp47VhE5
mW3O1Rm8kD0TnHBTiXffJPRbuOt05fTkmXe8B8XmDUpfWXLDjeHjWBZnTHsNafnXy0ptL3fH6qvW
QpAfu6GRbWRFYgGNNiaWa5mX1BUZ4HvgylhJS0xRJcOoY/vTAedXndIbLy0YwRwf0ovhyH93M8CI
mFcOXo8b/5MBK9fHXziOa6do42Vutx90LPr/LatTMvmGMNZns306MOswmkZaSFReXab0k3BE3tG3
jb/AnoKe5ofbwXKNAzlBLEHf3AxPjqFwjBLclv8U/ezciWhynrB6OyHmHxtp9yAGs6Yf0sqrqabo
skLvJts9SoyVx1a7Hwa3BQL1at9aEHzo/CL9iyidlFNKaB8ox0RYtzjVDKrf20DMIfmBGDb3VrKM
7fElSXituMLJlHo7ty1ty+PglGLiLvasCYMnAENUbtSL/kJVaYJWi4xeWgLec1GHYSMqvRat3DOf
g0IO+wr12UfBP3r7amYcBXUOROADWPY7ssgqQ48pDKnMxK7JhN4oI2Tam+RAAzXKD8LFjMiLmIvQ
EvvvQzH5Lw+XlqavCwqyhMiS9FvJbL8hB+SJGCTpiDCAlaGjMM9gy9ClRi6KXqPaWSRT97/mxiVt
bfQ4vzvV5gLBrAE7gZabuFp1eBCeYhqOT/cE7CwwB7VgTUaLWno/CiJPQKz6hSJOkT4Cx21YJpaU
CV4OdAZHlRUP1oz3mCGcBDAlmXJy6wvmFBzwnRUKj/McpfFThR8AcINdSu4hhEldmeNxxyqNK07o
gQuyuRKzATmeNpW74bM4OFT3L/hLEFBYJccQsYmom+qK/XDqqO7PXlbptfUaJ97/yCl9jGLHoZJv
sWrjI7B5S5KKtNzbEZnIP2U/5MRHAYoJQV6W5EbL6p2ZwjUmTu7IvrFyA78rkcbNgsyiH3atODAa
VDHHw9goJk/RzzfgbHRoHiP3OhGruV2EnTAN/RGyZ5ibQDLVUhT6GLt+h5l0iHx+oipKBBs9bJBm
LlRIJgP6JHkV7+WBE2xrmiI13QkWGik6Dhbw/vayAb8O3KXfBHgxVx36cUal5PZoA87UCqunl6CT
SQgVERbzKx26o2NxcjeKBvGGdjdd4xnrXOVRcfS5wopYZ0SDi7bgMFpUE2aAfANoSlIJGEmkGONK
1gvjjymxgUmHo7vzdsUEaaV9FgWsEiXLx2LSPb0+3dk1sMnLEkPJhxP19YuwgQU6LBUdX6DOLjCJ
9xIu/YEFZRn66NO5oX2MVBeQr08EnTACQeDLzojNgZpN/T3WEE8QU8TTPK+C/Yb/PoHfL+r3wVS2
8oeQP3jAgkrgCQLYQKWxLYbzsk360afbz+VREhvXLmckZIwthLYb/8Y1WzPff4pkRXkJZPMgTGqD
78ufChPYr3MiM0YQ3hqmZW+yFcXn8hsF0wcCId7l6GSswCq8YwDd8BWVsxF+70rnVQLG0HYDOLMh
H4ab1XqVqBa4Z3DNEGt4++08gCZHAM0b2ZQO90ds/6nx2iJR1JE51Vb80v+UcsN+JdXW0Ak7k2cE
QCtFUVFCxhUUebJs8Kifmn9kTyj2TQMy7Cb+mKiWw+DotGoJT3PmQ2+iIIJKOWiSEGe5hBZmNhzq
6dg5FeMBNl34qtN6uItGmHaybahCOiGURLIoQXna1/AmUyQr3/kfBI9IpBY/0ScTOeSJ7PQnl0YQ
iI358hI39Kv2TJbIoXyCqrG3MV/htfiQbddoxpkjQFx2OZmxrFVBvr/wPt0XNdwOzuJudMcglOBr
uD+tORf4/fXVchHQAIP6nHRE/6fbW7cmf3m5CEXfW8w9GTVZ+/HaRXaG342H4q0qStytJvZdVznm
Pi5B5rvLOWf5oIJXLmj09Kf4/UzoIgNSxZy5raL2SkL5RkYf4Z4TJySLSeadfYhF1tbgxwFZ8jNP
+ZWjAYNfL2LiMnec9zvJ9JclHaolWtsRbikj5JVuO+w4nB3TRIUoQjFV31hpSmMv6SaMi5ssmSDy
IwJssVoQONhsk8cT7cld4RM5fDWsgPKfmJve2QYhIOfskXWjTIgAG/d/VDxnWLxYOSVM/xbjzEW2
O4MuscZ5PomJJB+9tDi1I618Mz8yvYfM0P2wchAynEIvUxcgT8VIHyfanXl5z6y2wUstFxMvwdQW
P3S5YjigJZcwSfYBa8qSlW5eorEAOpWZijjCt2H8gw5qYJfgRdaLIAIbQbnUWLmyumH04uZ3nx48
ee3WpsAaRTUKqK/QWuAlm0dQs2h1MPH971alN4vwiWYdMEu/4E0KwjJ/pisSiOeXm0fMekI/EVXU
e1mn/a1e3UUAiD6q1KqH64Ebtic0RDPd7oQU7L6rG0T1fcUt4VMB++0iHd0rJJjXIdvJr7/FPMuh
2BTEC2MGy9P44Xft7+9XZ3GUL2O6SqImjB3Oz6moXww2ARwoZhXGJgEtvU3SY9fmmjA4OC59xbDj
b76rCcCp4iAzQ//O/uJ8d9JIug9wUnZvVQHdeqFQt7iPeWEXLeDO4dn+t+vJB+WQSn3cq1rg1BZE
w53wyJdrWL9zVsde5zvRPlH+POCJdb7NhNCYnfJH1qQ1t5Pd9GhQlffUV4LQuZvc08SdlQE2hWus
ipOhpd01FAhHToNQIZ04fiQRml30oHPYI6yOJksxgVBmIC+jU2UyQlTODzEKH8D325zZFldX2Acu
/NsX/3ZMEZtXsdTo0zkt8TJ3cMPJUXdaAngo6QNQju05J69VKsD/wk6VaeG9o3xTcAZO0DsNzrO+
NsbFqIhOLzUQvzBX1cMZHw7oHWBZgl6L8EOJ4nGbhHN5X+ZUKszoB9DM1CmBC+XQLshdXfi9W7GS
37X5Hpuvu3Pf0Z7xKbzy+LQW90Rk+tKqxRTBIzCFvN2gRJtDEKESFGmOQDWnRg4p/XvBdmK/g0Ud
A8kG7KrWnzBk9XSqRkwKqaqUeXBpTlO0m/2dLcs6WEbfNeeln/7Pfvh2ltnvbTWmsG48ZX/iq7fL
+9ByHuhIjWOiA3sPZY3g4isnRYKGfK4sqABLj8zR9wEygGrPPMm8OyXwWpzpk5yjyDHW4LKDo+Rn
+g7eLxKIkU1/RLlCV5gQH1Z28+08vWi3VsO0H5QGZy/EHViQzSVf3Fh5x9+UQvzfinpY9envoZEG
/X8Yln9Riq0x3K4Qoj3VL5yIznjOBUFtGJU6Xi5/ojeZkpOjTBsNZ0bU4k4SLU1NMVF3kGQtydme
yFKp6CwuwQr9TxKKh3DwiQ/o8LjCTx1BeTaCIv2108HrH4BR4A+Y5NYCPwwHVMVtjQQwxfe0F1EL
10n1MTVPmm3mcfyoM9jyDA8yKD9Tqq64V4Yw9cBjN6EtUwmK4luRGe9l3ag/a1NJUGrB0v6Rgnuf
tBJpVCrCUr7E21T2GFHRChP6oQHQbassRvxseLmCdIfP23gi0b/EkwkQrV7zxol0lGqH1aXbP8GH
nSs62TUYn4JAwe4KQ1TmJUHQdt1JsNiFjy1L026r6b1o6Yt+pjvSP72bv20xatSdKWFybK9/VhXK
JpjxE6VvZynhO4asxPgIf4poGpm+6U85J+yf8QUnt24QWoWlro1tg0K2Ypvq6FBECoXseagv3HeD
vci8Gw5kIJizADQIJzJvkAVPiyJCvWMERBpA4LkPFfbVbf9MFoTLvli+Oe166xtFAvQ4uOWCKfjG
iu8SeBeapMKFIdfTJzi0Y/TUdNx/6xT7smPNeeKb3HMIQm3A9W4zoQAMzRc05LwxXrb5G5s79oZC
ZSCBdWz2YTGSA+1zp+NJ1CanoNRQW3zJ5RGSxNVcXRF+Og/H+TcyPMxCUL7Ep5H6jfuKIJki/YcQ
dOcipIZYoLhsdZxfqxPMULOVN4dUeHPCrb4fAoQH8lCQLG5hW5L4yoCdWWoIvTK1I0BAtaNhBl/K
DR3qwMt+iI+2ZGl129mm3QgfBOEAeXl7u+7fhrK3LxaecIyOginoB5NRCwj+FzjEMna3vStgaK9r
9QjiWoMyqIDS35r6jS4zUdprSMTfPc7SF0R/7GpYTEv3h5nlKL3zexgKuJGq8/l0RajlMsik0SMT
/uvdE3ksErZZADnMyq/6Yy3K2JWf+YKzwZQNvI1A/nNc3d5N0RKgOlOaUQfwl8ZtkSvXm6W6Uh6C
MBTU9+YRK1ia8w+Hi8D78qHt49FstfHw5/CDxVlURmzjpmqy/zBPI+z8nNaK3U4f+oDqO/UcDw+3
+O+dTp9eW+/43+dpglEwgB8B8Tj228XGaUo1uKDGZVP2OmmaoQmQjQchhkQ8uTdR7jtc7U9Ssc3/
KWzTZKX5/O1zh08Ql8SVPCqd1oJgwoCycYYpwyHgpYE3xpiS2jk92oNWFDEGhXB0+0SZpQ/kmqm0
gSXXV0fQApGNYgT0g/SdsConYzvsxpNl2Sk42D2gGFVEtLQ11i4Qyf7QT+g3wB/WWYqtq0Tz3b6B
60BRuX+qU+fJnsgrujE79KiNW+8gJDTh6sddwreq63f/AINNyBynvUuuMIRvdHOSi6CT3ppJoyGi
mS8PokllS9SmklIqlfWcufJAKSYtdRMv91ovFZK8IDxtUA7l1xD+aXk7cI9HXBeHEc0ut7zaumxR
UPQDoHwoJjlK3uuj8GWsvlIGEGtQ0Xrn1G/BlcmvxU8/V4338yEDbezU3LwuGGBh4P4g3h1WlU6f
/3Mf5c3WTpTEOb/I/OXIf1PMr21tnTm2SiqatuSoIVnSrYdb/QU3QJ5ccPQX6hTh8WkcREwWdwnq
+zFWLAC6NJJhg2r5tA+1Md5W9SsT2+eiP10QH5QWiXRP755/fkbOmAuuzPDc5qiF+fIVTFGi6tBe
DtN9O8LtqCFK/iNMjqBoqezcz+G0fJDTbdpuRDhdx55h7hhrkY13/NWetf2SC4gpWbu6fdeRGSSO
p12YVAgF05Lv8YoUMZ8NPzKcChPRUUUJ8IY66pfQXv7xP1UzSdkuKBW4M1qwvDGKy6q6/fIDrC/y
YLRwOSduHLucIFy79OsF4rU7eg50uSXLhMW4yJUHmWN1dL9PJXDPfnZCMz1lc9B8qs8SBnP9EHA7
9J1cWiQJA49UR2LmdQckT1djExGaA/bxjNQs0ZX9BVCFUx9UOIwfCRIvkhO1LrNmD5HfwjJayAu5
6xozGmlCYfgiYBaZ6XQrSDTXCrJsADqQmHWhRSEUeOrejU6aYcBsIklYb67chmCH1phT9QuyYJ9W
jrCe7s7SD1E+1/3DwNx+IvmJrApMQ8YCikB9xIJs/HHaK0l8XWhAAZ48QnrYej1enbAX9zBg/Hfv
7yY5um+sZ1kxeHuUuPcPCm5kRF8D2ux8jJR/8kNGJb/ODRH9lHH/TltyImWR4XDtnOomz0V7zz5e
WVI0X4AtheCusxSxP4+9bbHbMxnNLdm/tW1ciNFy8T66eXDXgOwUKFVMG4OyBXw6RjEEZ2owVd/X
GfXEn/9KKCfX6T/A1Gw7VpKbYG9sB9PifBNqvVh1v48DUDIxN69uySijoDA9rGW+xuBHEalH2UDA
S4+hn1eTSgWOZgpGVPSsO+5Xj1gH9UCDVeUOERUBvrcvIOs84z2mjAbKKaETHn+AsXO1GaMp1x8s
ydeqR9kk+WhG4pAzffcIReZU8zYZlwGcf6xz7F8Me36qyKwoE/lmPDz66KhvsUOV7ZqDkTPRe5er
Te9awbG4lwhC8g43rWe5Uq3xkRnfLKQYWzDsLP9Zow0HBiNz/deLI1JuQ80xiBhtYjkJ96V611BF
II/3/Zskv1xPRfS4lQyzMlSEY/22S24cQOl73J3T6M0RY7r5mlUVCNvVofERj5fZCi/Hs5yR3sb5
y63FWb0l12xws19ZAW+fN5EiOMmOrwP2yw689BsLeeudPzJ73Iw2FAfvVSQ1HR3IcSXSRT+Es247
oGuAzf661J8UtkxNOgn/5lVsrELqRD1cBtV5HR4triM33KnkMe9wWErLKuuWuGPIMCOAv189Rvff
u7Z/G5QZvUbBIlEPKZ85TUmDOzTJxaSdawQhL8PzUkVWGXKfdj/dbj5xrb0aDQd2P8PRHd4mj4gn
PJU6f0MzEoMwZYZ1bOsUPM1poH3Ehu9Z0anWSzwwmItrdWDG7NIydRBj+WgZYvksK5TVp7dWZ7C3
XiiqE/Thg6thIaoZ9ZlxwKTlnR8y8mWGbNNrDiMyCajskJ292BIHDpE/rBLNt1GDhoAJbIiWbrRl
CofUQ72gZ6GezBDYNKn7RM4dboj17x4Hj5R4Dc/COuoYDgBw9dkHkZBzjsRFmZXML4ihdnAA6Zsg
CAoaCfnXN+65RPJaGcCBWFiY/hHknWY20GsslMQtUrjfyeTpNJ0LFnCKdVivFmpNPNulWInQQ574
dcs+Z3N+AIQNl89wr+IS0w/Ig1jXlZtKeD9emPV3s2GSojpFSlZpDKKaHtX+eFiBWQfIuiBN56ga
TXyVeeuHPDMDW0fW5NHgV9XqOlUOwwv/YTkzBi/FoGEz7/vXhveD6HUKR+Jj7iGrQlBubK/lxyFF
9hL9EckS7uNOdklDt4aRBLqsmxXAZlD6Te71h1NaZf3qbHlQ+H3DPJYqZZklDxj3hnaHpVsIRaZn
S2LTIGCYo+rhPmRy6O2E381tVNAyN1B/HkIVVBRAiY+TvHXjWAciTY+FV6hi3s2iH1EGTgE3MKvC
lXZwlKJE1NP9979LNLtYFlcLzEg/VqCzBUr/lOH4i7A0rARyia3rCMzx4315Ap4Lh+ilfaY+kiPs
/BmCS/N7uvyctC2sTAPxRqadAw2nR8HCDpQY8O+36NXgMpNh5I1MKQGrB3DJxOgrhM8FMnL59/ep
rHKkPU3czduyUexS6hCm4LTHr206jUQUZqGhnSb+WfOaIZhvZdsQyBzN6rKeGB3WXjXlIw7X7rZQ
mabJ9NeXs6fBOz7czr2IvHRmGstbIygIxFBXxfbfLj1N4jfZfky0nHk3vKqNXKUQ+8/kMIR6ITHp
kmY+Hpt57BGcuKyVyqDFOEYDYNw/rs3lAfzghDlQGyTSiCjGT+1g3SheKSpn0jkWZv5AHvZCBpd1
hzBu+Yqd9o4Krrxv6ltJ47h/ggXHHq7PZO123X36gqMiQJmqzRlsJMUWHqE8pfIIqM27Vw49AHAB
cpY4pfwqY3016zY5x8RwDBwUoP3pPZcCo5fezbeh810TXrmJCbLK7lUkoQ0G45Rs3udaMOEpoOTv
xKc5cPa2c/APofLxH79tR6sq6LvrZ848nGGOFs1RfPHzOKSQJMRUJy8w6kUSsvjc/nAIoefYUD0q
pZTvWbfJMKDgKsyIUxnpJ38wj07y+4nb2pJUz0F+v/sCs6/c4vXY1geaS394vL4kG234RSQs91d+
wn84RZUDseQsqx+g/Q1VuZQxksEm1mGtbx5QWkHUOlvxmGdhB/tpVH9M3k1Jku9F9XyYSAAKz0Ao
Ntu1gJNO4SNWR+hqzdkzngI126b4QJJxVl3ZbOyyiNqkh6tMW+Enpmp3TDqe3yLCNyh3W1Mt84QC
xRpJoO9slqd7X6V74ThQP7+vVQ1isPWXVoy0d/YctD9hI8+i7iTevmXZHSbrXAkapin6/+irnG9c
v0HN5h3Pdf4TSOYEmaj0ayTKWe0dEnUVzDg/yqG/cvshSQZ96bnhNw+1fvn9+wYfP4aZTs9+DsgA
ugWIiO4ZzjMaI/h6xrzcjCM5JvJU22QUd5qvNTdU7lWmANo9cJqelymEfOUefV15Mm1ArxwRqjwx
YPdcasNI4Ru1xTfBJDSJcaILL2ilwkjEMI9o0v8lDriod3QdvVy/4Hk1AyarxX+Na/TY3Ly940+Y
9sYIs242wp9OHkL2NyZwxGKJJuDwAuEqwVQOkNRITLa2N1GB4Plu4971DbeBhUhpiqYa6QqDGFNI
xVJgkJQoIeCDq2UFTeGxXkXl14L9gD9nh/qjkjSsRI6IrfYUQb1Gmdi1e5BRU64xDqabBupU9VYb
FYjNYBDmhirjvqadCvpbv9PYxCzBrcdWWFrrEThIjv4he7OIZF3650DqZhdsaRTEWp4J5u8wYcSe
dh/dXJUPPwSUwmH8HCM+jJumSiF5DDM69pre4IsWeUZcPm4h9WfO0erXEPOkELYJ3uS19NI4v3pm
zi7yVmtpwgknGWybwVSkpuTD8q6WdqXeCAATFRlq5xlnSZHPE6z6ONd8VIdZfYqZ3+i1YQlEFnqA
DaZaqXPMU4YQPPIzeLcfwiQDDVUZNUwZfmqCotqdoVjb1d9CqKljNNO6R/t9pGBP1M7/yAWCmKaD
1fVKfZXbwQPEgTIN5A4I8wchkse5aAOhlC5d0AnqBdTxWhtKtCkzckfmQMxLgJlROCMN0jeUYHAH
M2Blya2QuKHV7KrRJRQUbG+WlsTcFiay4rf0D4OSE32ET9mmc3rLBREiYQDb+FSMZF+ygL7N3HJp
aVoPc4awrZwbdgPSHU3pf3axHlhI+vBEDSJ+UfB4i6JwBegyf3WWKM90Ey5D9+GTmrCQrk90uoKZ
8NWDuJOkGnXl9dazWDWew+QGc6vJj1qaefbnZNwXi9OMEIL7Yznp4go1aH9Np6ibpiIXVXrxu4iG
tkhPP6GMg8NqGBgHPrXhWyiN9rqRCUuDzyGKcS0rbK1P8oH7HbWmoJ/k0RxPho5x6FCzg1TLoiRl
4o1R8SEvOKWaRch2ZDr8P1gVeijgQFY97mmlgwELlDTZnFAj111ni0OEP71M0Tc9aoPlgE/ZcLcS
qDvQhE2XAyYhaLlQ+Y3cYmT7L6oNpukjgLhMBtZQH2eviJ9pu2R59vUsMcBpL3ZzClmL2Ve1R6K/
RIDRURA+hLsIZPkK7462EIBl7L5DZ9el51GlK6NdCruLIiLYc5/OR7vLURNYDeXtwcgr1bx2bCym
FrysR7iFpD63feMM2o41rpBLLsdzkGa4+uFxb4Q7rIna72WGI2uHgdReeec03A264BFSv0Y4Lr+9
OD7C0OXSOqjZptdJl/9SnXLLdDTSU08BJcwoGuyGBQup01ff6NA+QhHG5TK1Eki9ja9wS1NU2U1K
niRjL1bMp6lebTnBg1jkElZwmlo/PYNqj0+zfr6a9D2UMh91Rhr+ocO9HFRhvupVfCiNHID1UO6h
m5e83SnqAmCEuE06sMn0pYqvfd+eXeriBBl2f36cD2XvLPZOTkZ3rEo3p75oK3QSmYs6atIpJFym
qaoiJN6ubI0DVayuvLXXuV4GacnZO9TXEnFm7FgECrWT8wyvmpv2xUPEViCYtQ7u/w1igFZeFNb4
J7+Yn/OLY9CTztUGHlPtRLLyySYnWNehcrJgzR7DHSzHVxBEHAJR8djhCeb58X+MyO/kPiZHj3Jv
VcodLRaUjzA3DZdBextR+YsqDQzKcOiSjExQqHy16YObxDC1iQC5thfhmWeMqXXQ74ME2LRY5XeJ
P2gAV0egaYaDUd5iokCx4Dohe5TtRV6t4ML6gW2lZktjBEJRYhPp5I9lYtlUHywFDfpVvCuRNBhW
6NbLOsjXJwXIyVtiTOsJAQ69BXSgYRK7N3OJz+ayTt2//86177uMrRmK/wITrbeK/aqrqrjI0+AR
h2hqgCpBXAFSnLALVryyzHRJ210at4Q5qZfSbJ3EpvN5B9RlYBVPOOtI35I6XngP096tSsdCGWrA
v1gHBCR+SYkPnR5d6BF58TmTre1GfK5bwWApuDqrj6IALgzDKRptbu3N4JLw6neUZtFio2I15Zl5
rgDMgiWQ5iRGXnPmLArX0ERSBCPURUYDzNIBxuvzHL8El5dJZpWKJsNAcB5FsuXoCvQaKxkjzt6o
Prk4fb8Tr4O81cYs0GuU5QycWYmKsTksvzacNdhdtpUf8tkzbi04penwSpCFkIvuJaFEdYHDGNPF
62YA+f8WI5YUBn37N46aynNRJ2Ql5EV6y/+ErCOwu5DG68i18f4TDBIPjaa1sUcr5JcMAylJtcaT
uCu+QcR9OGZ9KI8POhC7vYQg9Tdpcw5f67hRmpNP+6qyT7ryB4LazJACGs64+R+j7fSW27CW8VNZ
X+dcg3CM2lq0fgyk3SfeOdFKFjzbWJpOeMJS1Ifvj1UflVC45R8Yz69wvU5R2qLwYzplJzlxaSNZ
PzXAsO1Cp7JyXkXdp+jScXg6rDPw6RLUYtiz4BcbM1ZpnCL+YhPcA8qumiMR+1iZZhK0hcTD1kU5
m19oPrHPnBUQx4uEZ0Ra14jbFOvoDwqmF7HQ/UEukfcQZQB1zcfQJGjBFe2xpL2t29uYEuOLwbD4
mqNnOuQN1B+o3GUrHtbkG2W3h2+sInhaTPdc/xif4AGq2l8/xkGdEdtJy9pQWVwiPyRuoQpI4fcK
zvakEbuh9PmrJiiGvQB9/DZXKA5EsGzU54rFSNZ5gdBPxY+GlTvRUEmN34z3hrylCWsd7sIPfWLb
TxXLE5SfFb5dsWeLzlDKqwxU69g9teYsqKETivmPEa1qc+j7G4CjOzGeeMxSAJFpWOBACjTwLyFd
FoHVZte0kllB079q3bIlXCp4OVmQYMl6cBK79oyOfRMCjKlqrkbJuO6i2IYB1chHtpcKuAazZgwV
VGx1ccRk46O1YIm2FTNeIRyL6ISLW78nZOcH3CMoo2U7Fjn3SIjlfNzIVnx75lsIU6RBm1CSazcW
+W/LgBZFrRqBhLzOiOvT9omriYeXSdnL8EujhMJlYpJfNK2Z4pHeR6kS5z4RgZi0yORlunQ/sicj
yvFBCvj/8amZ1ZRwWVCdZjbuzykVQqfyJ+GJp5m43q2bVuBuVkYJLGLOsJGzUPKP8q3qmnxI6k2T
IQ+27GW8dNqWZ4BibBJW8M0y5F5QWembzKWJO452eyGkValSO1RdqDaL8mrF9+wxw91+N4hvGk3Q
0yloAJK7nrQMQIKgSx+7k9ysnaWRcCM53BynoxoTyp3v8sOLRCPbBeo+y0Za2Qo//a1NF1hd438b
uHKQ9xC6aD+FVXV7f+PSY3AYDiBSeIDR47qAmcnplL25gsaqVuWNe23sP83wmLiRfQAfvdle+IN9
WMvmVR8pNPXfHqR1q5Fj8zGgcTDbCI8X5TiocidLN1fNhdEEVj2QqmA7+RS3sEmTpKREtV5I4ipe
5Ji2aDt+weAlpXJhIrsn9abornNqiMjLu4N84PjJDQxgaisv6DYxQqyLJIVxI0cWRgOtfS0rL8K/
3uhM7VAsOwKh5dozX3L+V7inY3wjU5YqdY1kv07uKosd0kZ/HwcwCw764vAODuOARIseTEBiVE5/
qXofGWgmE797Jyfg8ugpht611yYAGfndo7u1+yQyHZ+Sl6fYWgzu+l6YXBQ/2okbEnux/qZeta/J
C2gbOGwULC6obV4zXtYkAlgrT0/ZuN3mUTD/TtPPhrj4ng7ykh7JB0WR3l8126xzYpllvzFvVTl5
g0V22odEyrvil1K2Mkc5RSTZMoaUGaRewt/qEgnP3Jg0qWZjwbViYd/59uMjeI1OOt4u/pUxosGq
CLQGDpGWU9Pip1a3M2Ymfv6E/HHoCp4WY42/savrJ1VbIJLkmH6+4m6QgXoEVIZ2OS8OcVntGqM0
RZbfheALbklHwYjrFsCDEfSgM1P+jAtQy2g0stgqpEP/i8F5UoFUp+3fMJE6+PM8KO8j6h/+6enz
X1WASDzXRGnZAIVgwdYE0IMpuv5IhMFvikgq30RVX5QMVM14N90OBq87atEaqhZ8kH6oBJa8EV5Z
MvFFfnbxOWbd/DPdOMMJvbe/WnVYPFNXO2rxPlZOJkA65Ydyl0FS1gFPVwGczH0+8rWgTmUZ3lbD
srx5UTyuSg3xT4m8ChlUfA2l6MtaLX9MrTjii/GQ4Qz6zLCloUC3I09Fkd8O3TXM6UbQvmPGNzmK
va6x0bWsVwR2rOw4JJt4ixDHKVm4rVLn0wJVWrXAXkpkJEhSHxUqvDY5++qdU+9jLEzekewacQRy
/z2eScSkx/Dda2tzSah3WwY7zxz59VtvTU5dSqVV04meJcwoGncQyHv9Q/QNOmoXsSAVYy2wuhQS
YICIotTl7bV9S9nsOs9FaUIcD5c2VAtJlDGXbjW7nAyeCesMOb7nHacvveupNVyRBzgRtlQcAVoe
7xtmeIvquGyzFb/f0LdKyRWE8pLgibjrlk77p2avzUxdDfHcbCdQoTLolbLEviaOdVMrXcK3bXc2
6UrZx+LWrLD3UQMW6IncZ9FwRzUzukHlOey3F7ADwCO2o16XN8Z94Z6OoqMSLy7qgwKG6G4c7fW3
UqqsfUUcw6NCNRr51yrhBfja7cp5BHMNSu2aWbof/qrWoFQNCHMFfJiURL9BIgRnMoe1PeVSZGth
5hHAdUsriBq6rYUejNNkdtDr/9L44V0rDlHPRHREETdhUT4y491zfST+4LsAcdyZ90Nojxm4YcYt
FQx7v/Di/92NOgo77O9vphTdq/d8DXXxonjvRMzGhahHg6Ngf273oPGHe8zABINyj+REdlMBBPHw
ljVD/3lFt8pSSxdxbOIUGOEBZAqAoGswBcbtXqBv6MfzotAqA62//Kkc6ILGjvQEG9+gA6xg60b5
sZn/T2E8rTsM+B1Gi74gPrhnJN/q0HLcA+iz28k/YLo4ptg6X65lf7l2ul0bVVACQ4/rXK0nUBA+
LNMJwwBCVAs6LwF0PApZp0y/HCgUxcRm4AllnjFyPCFDQm82tOoU34JZ6+i40Hk2IuzWXQjLV6oj
ePYOaZpVoBvYN2iMmBzWnpPNSojR0StLsVPEPSDltGONV2EHCSqTykBx59Ib7W3FSS95VWLCSya6
pbQj0fs5pbQvZRs3nWPW0xEF/oO/KJ6u0pBRgmlpNt60aVaQcS00Nf43q18C+YxsAxM/D59pw18o
0MLKHC5/s6zmF3TKZiCU8lZDUXX93n68uHrBu4+epUELEWXgWhafVPjMynPrI97AIDIIRywB4u1s
vaMKSms8SGUtRjwZ2w0FP86epMoAan96wfz6dhehThDjXdkrNVFD0sDjQXTmiwodn9DtXenByo65
3oHfEuYutdpvgj5OLUZJ2UJYnLZW8QFoTgjg52ewgkpdZ9NYhBN6skBKVOElimUnHsBMTHg7KX07
QvXQhcFznCIS53UR4Cyi+ZDR4Gnq7TBsXjuPOjgdXVvolXpEN5bft1XHvz3F8qxApxCA6kjMlcWa
QxqBK98/sr3rY3zMkwfc39gGgZ5WJOPpP1w2XA5HLMrAT0hbXX7XbwjxXHYe/DyliiiEdH0Ql59U
88MX5zWj3EPC6jlXc/KLd80Hq189bel8px+ntz4vknFkXBrfEr4relLzZr8Jlm9IgqHHD789tIoc
hRJE7AjwHX8k45nkwSNeRMeMfvcuvawgpap+AIE/I1Ysdw7nLVTcg1/mTssqWHM6thB6HvHWKPWz
FkMgr02WsZtxuCPL2fnFPaBQG6YqVkgVj0OChcseRA0jXy31x+jAoQodhboAHpMcB0zLioA6B8OU
G+4XOS7Ms9vb5j6eLU9reK5pWo0RZOWK88NXx7tjwJSqbd2JK16qVprpubsTJFyGje2N1UYNwCxg
lKVA0ztDHiybIwxo3QBUmMr6RVFZS6GqBz6dEXB2/FWIliVrtjPP1rfXq+XWBB9f1GB+6TtjWvIg
Xq2XAiY2yw9Ty4q5NgVSf7mesynydouDdQWhuX21YdKbShOiu18/sM5Uq6HIyMwVv+S13Nj3vz4O
3sKpGYZyPpN6/ukRqArr9YQE9pRNj0PaGllBvFKZ3zntIOmHtxtN+xgda9P01n2YheMIYaY8ERAA
99GnEvDZxKZrwDn6ZS14EqXCoxKKDF+qjCJjWxuZ34SAp1+wJ0gF4z6A8WR/YmtJdh/5FB+EPJMc
GEQCVEZk3cQpROUCpU/d5bN5zLW96tbjTuyeqr/50EsMBz4OhzLbbyBnAF8OChzqIvMt6G1U+uvC
fEqyF7BNBgKBT0QxeIf1rlIVKC2bPw2ZmITu+73bqN4eD6wc+zGCDlYwp/DpHxs2hXwRHo4A98Vz
FhCkJZTFrd1DYerwtMCF59/aBQ9syuKHsH9yLO7unG6QyssUPa/cQr6eo1J0lsPKCYRdwxZIljV/
Lbob0USFPuPoWh8tMsB4DBQWKFZ9MAAW5GJMUF2Y0hSPVwR1y3CFTgOfHgSWpzYG5OKT6DnL1rfK
i8BXD5rjiZbbj5w4KXaMJUT2iVeiCcIwxG99FAJDkTyPq85vnBcTTZSPWdSbn26cXTq0OCMadR8w
XECUuGPgKfVymrlodhAmy50sPlVl1+7DEdpuU4cij7f+XTXUxEvc6JhueuGAWn7y7Uy44GFp4Edm
2PYeMfTIsFZ6NXo5sh10UMOR+DoxKXIVGw6Ku07YzjTiLEE5rtAreh63B0o0uwIhNafGDamGm81K
PGE+P4XbEe0YUXWySRn7Gk+YiL9ahKF5r8tSPq/krJU59ihEzVwJx9zOfTb1OjeEKsXbLdyHrMbE
+xwLjT9BUD8oQW7PM+jAkLV3roU+sYv2FvhinjrTXTgX01StFpsEr/ahVURL3aDXVas8SiaCdfBI
TdXV6VCdb3exlpMA6+lbUPjUhOl49xGIvWXYeS0A3FYhm9mgExgIBsnY8xEh0YA1gBnTx1Ze+mD9
uYNc8TRnfpd+t2AKzF+JTe0rggZmYdai/LJXFhD1kF3oK0Srs1PWrbprWSrrnkJdcgyvA7nm2zLG
/4lPKn1PE6ytZfXahxgYsDgxqqf6/3rI9eBNV8EwKccb3Ki04b+EsblyexLHC5oe/oMPyCyyCjvA
FsJG6+mo0mAeUQEmvLM4JVlhKsVji+x4JDslzs8qd8IBqCGDU+ztWj1FUgAAeISxmd0LcPZiX0jA
Gqg9Z00ayPN0dlwu8BiiVJyWbxLSxi7hryyczBI+aKyxuHatQozD7gr0Ay9sA83kHRpJdjjhvc53
dKvxh7C1yUayVNKyLTrznlTOwLRCmgi2HtP6oeljjFuC0IWi1TCHVO11y5lAH2wrCj5tBcnEUV1E
npFtJWkiTncsoC72d5hJYMB/urPwmzKPh1Uj7mBAzlEgw8rzeRwjHxyWFarRWnKiq8ikiuu0fjTg
TO1ZGL85VA71soL+lYuwDghjq8F+z7X+fAonD9YsYY2OR3nYzmjm8EhuCOnY0Aut9+lcq05T9/By
qusSHVLgRfW01RRCL5o4uk+FVIsd8MsrJ8zmInb/18yd07yFh4cUhLC2PAsEA+JroggwT5wjZEfy
2bVYqvaIa8JtEEhPn8LmwvXHFximLY+31wd1YBkN416LXmK6e7HsjTCiS8BRf3ULC4RBQjxRzVSL
xQlYMct/iSWvj99X6wiYWM3LvY0OsawACHOtexqWJ1htQy2+R1B5sWAPigxLiFkD+MgkO5DtigfJ
ERRm230PTRCpedJm33PYN3FRPEwi+G8g14Vx1OGlbjV4ulG6rP6kWjuhwNe3LAjemdTZKVyGua+6
RgdpqiFnrf4tzpxT5jTWiKe32er/JaN38Vg2wIp5bjkalOnWtt3DGvg/OxNkft+hQeNzpNPSgSbh
GrV8S7Tl2CxmY+mfruD9VvGOSSsmEDAWszyi3W+CVRinhinRQBzWalxZO5vL/DOV4d10XBYUQBfB
FP5g2JtQKpIkToDpNT3O2qFjfET1/stphc2Pnv5NXAvKbgN226kNr3DrfIurJNdffNszYCfX5Ttw
BBFDJhqvfGGcidHaxf+Ul66nyaCGuoode6jrvzatmDhCl3QRk4HRlvVMJpyFWIH3wH2UrE/ad91u
z898CiXuPLPyA9MZKqnchkKCzz4gN38yMPVqDquuJ4F3LDiUuNmFz/QEn0jqwx01dPPH1FEWqh+4
NxIt+BC+XmnoV99EE7+3XmRfnoIwDj4nvDJbqZxtZ9Yyv7v2ws0OFiEnjC0B4QGQE9QI2YjEk7vW
hhxXNf5BI5jWbizWzh/fI11oDEFtaqV6lnt5pXBL1JGAH1fdc9sCJLMZSXhuUHQJCC7a3nSwwk7M
lpbD1wQNiBkBjDjYQR8NGIYEtJF7Wd/ufTYuNrBXTSx9lhqYL4lCDtuwHipfxdnf/k9Gz9aie9MC
gtyiX+qNzKAONXdGjl6ZSdB30K85Zy7X7fTzK8uNLQG7rq5OCOrVS71Q8rx88+u+o6AB2Aa6iETs
ljhMovgCn3K4U3eGiX52oSGJ8DcoF7tNUDqOahEbwQM9Cjk4zykzIpgwHkRNv75FT52Co953rPi1
yTX/2KR7NxjjQ56e7fGeMrKaxOH8csg81wMxTuSsAB8ID/4LHbQWr+WsnCGJi6WtI9d/Mun2tb+9
JLVTOhzfTID5WoZI8QSUH8fNa8c2+AI5QcxqoSs5Orjggq8lu2vQ/UtYS1OyFPRAd5eUYxPXh+5t
Vmk3rdFB7UZ5ilQKLpgZdM03C1+iHwSlUxEPGwyvBAceim1xXzY+/p7NszuEeTYmA3+RIPzcCYwa
02nVyemZiJsA6e44B18BrB0sfw86j2CozKiy3iU87W7EdB+iq0ltUcVzPBF4/uZbcPnP5Fq5sCiP
dwDhlES87ZtwKyuFWfkysAbteEcGOO2iyOejGxUeBP9snYhaxgLo+9EvKRMSNeVWlSbpTP81RMvh
OuL7lUkzhS6An51IF9Z0wBZdpq07N7xIc4VPKRX/vMRFg6off33emejBvbIMrOe/KPf0f1S99Fqs
kFBTl8X6c0DEnlYyUoZNf+guRYqePtVM6+2p+/wA9qnrOxWRTA14Kh9Vw3X7g5haCarq6rUltM72
mFNle57ORkwjtb+jSjAC5mHXm5WRJDZPvoqlPVCHEurzr7OTOte1yqS5/hMYui33fCTDJGvaWRfu
NRM21iHgwC/dQ9I8QGIcIyF75rVYJawDVpx4ztB58bsQtopFipEvY2B9BE8mLhKNFJNRezDRWONX
e1H12csWQ5JeK7fOh4IS4mDjRkokhHpmHZGQdf7h0vqBFRQK+UQt9AsQzkZL9ypkyDIiKIzdA9JG
/ZKm+fMcpeq+DZbcNumqz7URn8YIUg8O1XYaXQpOahL3slZctLF2PKgyuJ1b9ZD5TdYevGxrtvl1
Oe5HfLz6zH8G2r4Go1N8k5gxUlQ7T4omQiITx8fzAbX9NcviWR8wZ4L7lGTtVshCaivNA1Ft8muy
ouIXW0wdAcRkdCR3DOxkFIxmsa25XP2zU7gJ0FtOTaXCSLWrkWLz8trKQuiAjSluc/+OPRuyIF86
KECXdc5pGkyohz5ME+HFG/nbJLwIquj8Tvupkay57sRWJfGJK3HlOz9Yjf0uH01CKo298eSOsFaY
1isOsd+SaMndXMtlRxZULhVDT4B166YsRXDs0+h5KEdq/uqIG+o+6USlIHQ+TkBtRf3XO88/bMm0
adtS0F3khxhdAP/QsJo1YAY8XaWp79ZdckVRN+OMiRL6cvbhRaWRT50i/vBUkBF/tThvpge8i4gx
Pdh0UG5XZ4LRACNbHAfvJO+at8OXO+7EECWsztz6KnXszaC090YfTM7zMZlIQyFjV7EvM8W+cmuz
9529sR0bhceadrlfdMOfEnwOl+JSbLVva+C0Z4qBPzhm8MVTsg1Fmi/jJNb48kHdE1hoX1VO6MjR
njwNjWEVtAGr7QM+2nf8otRjXNcNAs2DSnn+XXCtSUlQ+QkrOO6vuv1xDOYBzJVnG+9m3fCT9X1D
wL+fCUAVSY6EshR+B5EMh89kY83IOHjOY9nG6of4BBMi+Cd5ZYjwwZbr9c15vVeUyvJzyF//5xjn
pA67njNw2A040MSAbcSlM7Y8antI6HUvma4C8TJOFiOX+emtop/5URXnsQq25PqtLBtaJT77Qx4M
aO5zA/b9FAJORKXC+Tb7Vew3vfhi4CdQarbrUecbNqBzYX4rlZpmJyUNckBHALp3INESo/QstwGu
wcH6+1cCHAcHPQbU4XpmHKbbd9UYSsx8tm/FeuTYAplr7bPGDHU6cJlj9IJASpHtM9sQSU37z3pu
BDpgoPsJHBQGv6YIzCJsk74H8SistU3xON4NvH/dfkqj8Xamsyf4bET0B07NaEUv/mq6j6/VqNe8
bUrVmgG8o0rMvSPY1s/CDhI3T4wliCH2Q4+phM94iNRchjhd4H8+B/7D46zeA0XjnkjTRbP+djmN
/55ZsFKu+9ZcwsSkKp7loI4c2ww8/vCqaLV+uYy1gbmgNotv4TcW6sGhDetVBK/Wr6uLOOyY1Jlj
gdbAIqd/ihPqgewdQI/z8d30RETmgrv9HQUk9jtXf3g2F52IaCq0OwsYevYXG92xVHNgCLwsDW4t
NZFZC7vFPFmY08+mZRj7imNggPX3/6Ed99ea5xFHS35jh9ohPGzOZfhC/QyS39RmgXXUZfMU7nnG
Jcu2jHHJpXBtgWMU43T2aWwnB5I68lTMKzLVfdNTuzgg5PkFmU7o/eTYumkVLKeXjd8XzZUZr6Yi
YnBbLwBdIaUwSgrjyqTE/sIPR6GYKWSZ6EUT9MY+3BPwcDLJxRMNwDtQhJGBMY4lQPHlbRREz3B3
6R+r8rEsnqcaEFLvS63iTjLhhSvw5VQxu+B/O+EJImCfSG2KhH4k7GC+Ov0Vrr+eWIJBTSQolULf
nABfJVFpYCSkJtVe1iVXa4nOZ134FweZzyhOOOVUSOUZvkkrxkCTcLacfc5aEoEO37yUY0dLmxHw
2zWEHekuhfqQAmfMsB1+BGNDKF7EVsq8H7XD6JFVkfC9KnLejgWUhPPLMX3j/pKCpV9yiUBHVfOK
p7t06P/e5puzfSBzcgRedJVgGhYfulPFjo+/6THtatemkE7O9Vj6gPeZFv/aeJNjfl9GogW6jaQ8
UGdl2OiRgkdb7ys5TKedGAEVFyQr2JZj8PyR0VblHt22elzxYdZF+3pzhSPqXDW5fLbYaxXwrSfq
dXZd5M80J0BsYFiLWC7gWOSzFAsQ0wJNpLF3lBod/U53qomXjWlbxv42sXbBVa+HiYJr3XTf/lPe
iejhka+Iiwyj/MoC1JZEZUR4HSLLGf0pG/+oTATXMFX/Ksl6nzwpb8ChPFF1j7P0J2ysg7aPCTv2
QLArpu55iT8sDDa1DA//PmJDoA/eNLJIO9XBJpNLbyKPofDC34XzlvDhGtFhE1qTeV8TELKSmIMJ
ovP8WELusE3o5Q/fiIxIUXSzOxjIyK9O3AfxBkzpNeAxsAm0ExP1HgIfDWLtkGT7g50bX+Rtipb/
eAAnxGWGMlPSfNngkeEmAaxuumJtOR4txpg07zoQx1gRgtBLVY7xMUhy97wS87+fS+a0IMjcaSnI
9peMgLirgg53MNVoSoC7QfhTmZaz6B8IVPP+Qb8yPkc3IaPzONQkUQnbowCcYuQlPkKANGRQ+2ZY
N6U/hW+9vZnTeC558Ze/EMIi5cOQxbPg43ht8FQUDtB29UXE8QGkT2UhJvTGjShIwq6zjCk9smpG
p/GiEB3j7FDQ7YAfthp/QDeAKSpdvQ7Ovqk5HzKrMZbXn76gAmjrUxNHlL5tHXGITo+EOsJy/yQo
Jvq5XXP9HID9hPVEemQrRLPxKC82oiTYCNTSAtgygg9GjqFxNmQAghwJzjmmbbdnV8oNUTjXnueD
byZkDdkcT1VRvpZs4dP0PMllx6we2bVzmXmSM2LO8hccnjseNa3MV9GrSa062XCiEjRSLvkToVFz
tQOOqYx5wXI9t+EVCqI8gpbaWUIP/SpcfIXUGmM6766CmSYObfMs8MpVJi6+tFE1/hippJ6iLRUr
1iMVYwWhgGHAECi67QKe9249P/9f5j5u7sECbZJGB+PY6a6ACEar+LCc63gwwHnhrEWlCNWqDmuS
1gPfc1qf4h4Xdt4fcGJiCrscpSgPsMo4d5D55Py2JUqa5OuwAJlWD7u1hbU1LoxHtI9t4EP8JSKC
X7mXhCAVJ4gMqOoFJ6Czca5uDApiOGwjsnb+VbjZQF0/VyDz0YPIyrdK049G8SlvEPCAuL1q3xWa
tcf+pIQFe+HN2ZeevB9w5KzTFPc9pwmkePEThdIWyfM13D1098AUBZBkmoYho63RrDrtTewRvCil
buWvelPTs0AIMysF3C8qMI9H0LtNlrCNgkaJR9Pdv/DLy67ZZGNxIU7BkhHkskNG7bIs/D4L8vhX
GbCO0rMo3766Lnq9bsvT+ABeTC2rwyHzS6GmRcXbfqykKp/ltVpzdC1UxLz2FEjFGbfcnx+iqt+v
xJqnH3SwReYKYt++9v2Wc+nvKNkDeHnFnL6ZuSUi8GiojabV6q3LFc2UDxlchMUaZwQgQlIA992K
Txm4Mboe0EYYgTJOMtZqsW+Uq1C3hFCw38tq8OCjXEDOIht5ZwEvmciooRqfdIpm8SO/JrSAodPS
mPsUFT1ktQoU35c0olH9MsYbrc25rkA2KJpqz6VZpYNvNlhMRJfHYl1425VMkkyRz/h4OVA2ob+3
NeMysxs6e+8Lq47WuSTdePaqa1pyhadBwPwX6drGt3oy3xSvhhSJAY/oSuIoRqDC4slpNtuQbArM
44kQ3PWe4JYg3xgBYDl7/a74ieoP70rZHLS7B4EaK1HRW9g5WDGH4jTh5mnbL6f3pZK90hD1oNso
1PI7uuzKsGHFbSpogmOqticeqJy8AepjCMjYNaT7Ta3IPKgSsbclrdJCcAXC7lnKf3aSzMyn0AWa
IeiQCLkikRIsD3gIyaCUvcMXMofO0AJsIua+Mf/IP0gh9DRi/Xt9UYTzakhLuE8FAM39ZQP5maqG
OJp0+Ydho2OhUTlY/8a07HKZGiMWTaBQMZV0snYCy60TRuVe4QaW1nsQyhUhARZm9/um2qbGED/W
oZQJG+6ebcVyN7uI96BcDc+rWNM5aD60yQzayu0FklElxv4eyKmxWkXNlBrEpguapWkWGFOJNvJZ
Odaz0VyNDssDGYQDcP0mBejajcLUWFA2ITt1nkjx5HOTL6CAxi2FEf7en/eJURwPcKlpTmqveno9
qO67rj8R5anaDMO42m7k2qwA4KJTGAH2JxCStPsHZnsxMiOQ7Yk9tcCXnwpVbzubGpw7OvgwpHGh
CLKHa/T9P/0MPjJiMMsvCxUKidGgDWfJR3BouPTMlgY5hqQfZZ7gZXg9NGET3hHi5PB4Gpiqs+wK
eFm2drn5mtty9IJ4FnYMonOnfnOZs4CeSjbZoL6i6Hq7FSJqETWEMFbu1q4HiQ9ZqNeo/37Dqbq9
RKvV7sssJTJkE4/ik7OZWCBgcF4bwWRu/2yV8Rp7YQbxkTRcQYdLn1wDl+Ug2MCY0Mh0AlrpkKJj
xDN1aXW7MnXEE4ljd65lShpxJWL1jzD68TbJ/Es52rqMEm8wImgnRAH4vxHUdd07mfjRO1nhNxAh
gv6R9ZO9UabG6GqufJw30ztvw9KiucL7fMtKpGSqJ1FydG4fuKXIgxH5BXOhpu1hkU7dcW7zzI7W
fUW69dJif4k8bJlm0kOZsPJ+/fDM+9eVm6MoXHjvWWJG3pkQgZaDlRYd8bn3flo2A1mlwKpMZDN7
Wcn5dJKsrOdJMhr6lpw2p+K9Fr/QceRpMi8FtG1u2GwU3sOX2xO3//rcK9sI5Exbv1/RSkpzyN6v
7xtRdMBI8R+XuOY28fPQeZ6mnTUv0O1j1irkMFvDfeNv1hjI9MRQ38qa9Gk/+ZcaW4KV4ZMHsQQ7
pN0HBrmf+b5GZQS0y/NI9vzZWPWkOeUp16qQmI0h9WL98F64AgVCFyI6SqYM8c3vAGK0tAnhijRS
HiJniBFhRYEWsz3UR+R+TnbXfLwV6ymdlqAW/7rJssX9UPdUObc4s06tah6rQZDiZw++bsz0T96K
Wmx/d0hz65XZAlm4lCqkZTN7L+4dDJSi7DcuM0mHL5CK4jlO2lwjax5LltdXXJj2PF7PCZIX5vc0
iWmkzeWeMXNlEjZDVC17dw5rw4cLXCL8R92xQLKjCcAkTxDsLbvjZ7RKaxx+QN97v8GH5NAJST7e
hAJFGGd7Ek3Cvvw0ZDhnDJ4SKwScJpRNxQMk+6rBsqhEwXdaCgJJXDBxrTApwizLCJdAiMDE1bx7
Jf7z7VSQoO600W/tLaKk71zXGXFEspRsBDvWYkemoMZFbzGD6RvjErot7pxLuCXvU5Z4wsdn+lye
SQmnIaHl+KomATLpI6Qe8rLKPiaPAtFBZ6F6CdwEamHAMLyklqJEcV5wIzoav/mEp/NV+zIeB8Hh
K5ifOKTonveIKMOtjOYNVpwsj2sdBWVv/ppzeYWLilZo/HqbLeFr+qdpGfKbUJlOiG6IVy3d5K7s
URWM7LQAYB1np5syUyTZchOAAHBNzCD3XG4v5dCewf4mxl6CjeO1AtueWwTEHm8CVNBjh/Bwtp6a
FyJLFEMVOLTachCNuivG78J0Xhghnq+n0nIx2D24AAGgV3qFo/0oDlZMzVnBsxAMN/AupL3ZxcaI
PmvZNMg0ag+utwa1eoclmxn4vINKMoIii2kgzPL52cnSFsiPhECFSW6WsGfYMnyho+S5YyI9hgHU
s04arPAyVGfFctw9IvyAoLD/3IqGDOUYs74k6pmSGiXNIt+YQPkQDD+2g9zqvnio4va4qftYPRRu
QDXKoeiUnwdgDckLabWiXgiDE5dqy3udHFhTknqyVuxvsl3CjKPyOM7HOeFlYyOVRh+XFeTdCm1c
qAgBEXjpSzcjOEomI2ZXbuC5Ex+3tYUBm2fd74V/zTZWYfZhg216roKyn6NVc0X/lOEunQOAyxhD
H7r1zXtav+U3oFRt+l7KfIcAzThakud9QFPtuV2tE3jIAKkT2hZEsZjdV3aRiBCSoMfM15XHyM4M
pv2EKv4klETdCC2WmnPdW/pqR0yKxEF/GzO1aIuCw0vety6fEHDgxZU/VmESyDzSKIeuBevOWS6i
gr6QSTNQ9+1fWQRI6HTlYI0pxGUvt0obblRVrroQ+2bqVgB9rkjcsHlR8pjb/tEnfYIe5RcLQHTI
qW8XcikD34QA4G0viIrNlzMs0Y+DcuUh1uKuJQg8WkWGtzJucFvmdN8a6p5p5wVcUaGBcrpM31hD
NN4pFDcdjg+Q+NaTHlla96SG2Wah4dXDCkVNwXrmBQlORVZaerjsl8JtfeI4oUyoKoGrQ8Q1W/wf
BKolyyiL9AohR5pwu2q1x4hexcqY89rzmk1ntbWrhtbl2fcH/kPkKOQtgTJph5PF1E+a8yQRe8PQ
v1fmEyuK6vhyuXCGvNn02Sank2yzmzxM0Hh87xW8RHYH801t6KC7VPd/4jXHUk27en3d7p79aaec
2UgSQ8dHLjeGZA3xciKE5uUxUHSlahBUPEKxdiBGq0F2sJl0uONnLW2qe2jltlohdlcyoSfdNa2m
/QhbPiv/Y0PVdNoB2jzqkTby8ZvA/1fkYiPwsrX+732AdPdNRNb43JDTdcLbq+QGaias8uZAkJa5
iSp/mDf01Ie7q9U79ukvuk4NBuepMMMdGPkJGVvX1028M6QrAh3mGt+zdBqb3JGTJV2IjAdZoMrV
17A8OHvbT1Oqja20sVCISt3t1sv9e0caNrQtNuqm9iS4dGalRoJ1gBPv9p9CcYuODA6bz6zHg0so
fL6hJykJ/orbd5GF2ylhvTt+khaiOsrThjxLNcgo/CrtExXnXHCE6iLArx09vMiFru6nrH0Jv/VW
l8Ot50EDcvKUfRuryfqOX0nf5lMohktoyQ/0rySmLUH7vIm098xLEM9zI/I9Mprjcs4e4eOkW+k6
aVWls+JusdaTcTiNiD2D9tfeD50VX23zz2ou17zpbuajHy8tP8F1XPrxV1j7ZeKD6mQuXRpBS5ta
fpcQmgLd8LQE87cqO4wFefZmZHhdXHiOIB7MF1fIsQm0G6ydWltTyaqR2OM9kohpKW8wLPtGlL3S
64rYyohBag/7VLJlWHcjTShfhF/HK5IX+tuOhkSQMuz6qkVt+STnEQZTd4axg0owZlUPWj5odC6x
EpWE6nYlEev3Wo3s/ITDHixA85Q+9R+yddFpXfaQiqYDmtlC+qUeLDgqzWV0nr/qCvQgrWrwTwje
YQ7r/M7IuAOh/+Sw4fgtinnjpDJFjA0Rok5dzvbk7yUjlQ1ry462NhOXrL6LsA1hVKZXx1emvTaT
LOKj/kQAixY5vFoP2F/IIGM+BkN9xzGpZdyX2r4wSByABA/NDw7FOGhrfZyithhi1+2Jg6xF8RIm
9+y+1V7FaLV6hdtbS26IY/AmF2zQZcPfqwxLS8lAtYC+dkRnpWiGlvhwbk7cxb/I2O9HsRyI1IqU
H9wTixcxiYRz1FZpTjLSdLeC5vQ7pB0N2Lfvt176V5s8Nzl15xiK9W9jpaDCiaxAIhxhkxb89ZCR
S56eaT3TgrEntQyXX84xuKuzRCMyB1JnKq87rtlUHK7Tbu9WHLVmpveSMNabALMi1iezUmws4uA2
alJiwjz/zOHxppDSSD5ZgS1OAYKCPten6V3FBeigX3gtGNhSbu6fFsga2n9MCTuOOM5juaYRgUaO
CSjN66KNA6XXXUDPIJOF+peL+xyfEqwvxJU9N11Vx6loUM+GecTGmoDwVSVvU7MFTKy5hvnBA6/J
FEF2gWcYpJ8vZJ52lf/OQnZzbbdoy6CP+LzoDsRxr2ae9VRY88sI6x4+G5XvFOlmd+FT5dGtfGHV
V9kO1+oaGCib5ZYRANSlktnwlKUc8s6KfJ/UxF7KxGQNkvcgKQBrdApd11DjZuQrZRml0fxs5DzR
/UfYr3mKXO7/hs93hbzcMGiCNo9NNy37ibZsBroFspeB6HjYc2o5zETJVcYx5KsxV51FHQzipra2
7Cc50s+/9ZxDuQwKzDCXajnsiFEaDXNQXsDXb2BnZ/5ATSxlbqdXK5OIQvMdcYGAqIOU0Eth5Nsl
+2s4phoMdu7SyWp00EmXfO1PqO642X9dOqJahddAYxyOyoMOmXB3fCwYlM6pMX353t6sukqO430l
1n6SZTxdlRPo+AVl7YmWAQbZbAc0yS9Z96JRUjbHZAWbGy8zc4nZQ5WprdezKGGT7iHruRBhEXbB
oCAoF/PDarXjCYXyGRvZv9wVq/pMPLxY7/W8+73epbRC/0okxChx+2tP7T+xTjrQhN1lGAInQRY2
HqnTI0DkIR3moEsMN1wcI6wsjFdJZFKvw3edRAA3noBxyuVx/Cf/pw7v7gD2e2SwsYE5NlD0tU0W
rwwmWwGhZF/6/jlg55zM0rd0vxmvYx+awtcvdopugYGzoG3yIVP5QWaxJIl8NpsyppTg7EBjnBD5
4XGJo3YPrZ7tPcfvoBwUpj/dmLL27BgC9xztIrFbnA+HRD9JGx6Z+AzWlCLNAvvQSgw4+az9zm7U
wqkn1MDDF4puye3dgF4EFS6QYF5ma0u0fx4RbFPUfomxSS2zspUw5Ied0URl/t8M53Rbn8H6uYIC
wDwR0K3Q7trZZ1jTkcPbKNU+sIV+gPl4HLinIAyohDT8ukv52rtOJHJktOGY62rk/lxD2dK9i5P6
/VFswa+QPFKTO5oAwEgf1yfxI16jM3ZK3lqqlSNzMWOblPPQM9gZ4xb+Sre6dkJa4HHeqVnxSr7E
Y2DVkSvz6MK06nWAZ2ZfY4mcJsgo5N5Lm3nAaXapwQV028wpgaaDfPdO74K5Hw7pI0eCTj6sDlPE
Id5jCEawyXv4uglIkTh4yOkf0zUm/blb1ltjuUFmdfmnMMlzpsW4rb2Q958iCscYWgHW4Mt22/w7
6g1Elg+jyNrHMAFpC4JC2dHuWDZTiQ7jsZiWaWT7vYGhpFvjzaMzGDRNyNVngIWcxNvV1NNFiDV5
46J8A+9v8gtqQb6sy3VpTI1++fG3njX/sSri2hNT6UsnBT9XVJB9HS8VXMZ5mFGHrltYza41P9Sj
ftZE+gdLfGWCZhIYvYT+PQigCCv0BkO6Wkir8PVw0wQe5fbuJ0yz5nZzXRXsXvs68t6zPGdd+Sgu
Vko3x34zzhwKqbVld64ANo+ULLZ4762ELq6wdOYhXsWXXcIcDeOE1BQpyIUvyQZApnD+AWraGsfs
ENydkH/1l4LcjN4V5GXkOUt5V8FfBtA9sNCX7wzmDMPgdx6zLYvV9g5Z6r0qLI3xMn9nyCpNBmjw
g4CC5t3qt85emSWyq0HnC+MIbavzmmmR7/nyJpshnY4e8zgSUr0CJRkpWXxcmFQHd3Yg8gNIJ3It
5ReNRsY2ZReSF9m9pYtKIKr9Fdtx5BfDAuiisWvgOs2ArOtiEW5wWoc/x1BlUCG/DGGZj6qTjVlR
2ZHFbZ9MfMFqp63YK9ShyToVSlh+cPftYWkkEgC4zrFWyNSAH6ZxY+1dulMgix4XS6gNyS2QzYwe
lq+gskSJwRiclCxJRjlN0WmQgQ1YgvqaV8jyHHIxVzl7CKinoixXPi7Ci2o9QBchX3QU2lx5smd6
+rBDie8bzXgEJHlhjkUl2+s8fGpRg/VEjWgfE8Ay9xlJcw4vVVkBEAs9ePoU8t02wAbvMHS6GEhM
q90oB7vdvHpoKet3rNOCethAQ7K25ni3mXBum4R42ZhAXLuE3s+Hta21kDAVnxSyx2ZLkaiMpIf9
JmlMme3yUHe83jJgtPPa2JRBONc/Owy43yV7d0jhE5PCC2awzJEB191q6NuChnu6fwZil0qC38ba
Lov23f1jlMUboHLIBgEKK1hwl2W+kTVW2r78yMef1m1/NpHBkzOVVUyGi+RjKzZBJZhsQVkHcIOy
8+90FLPsFRd2Sndwm2IPW5vmsGNHwmUSEkpL+GrbI9JlblfKqxGTxcUGc6lVRmNM9WQg9bL9x6wG
+C08CBkUOBCPCCyGGLQenIQ3ZgqEcFUW7f3zSEIKJZ1tCtrOZgdsCHlX8/J9/OoBXCUT2FqjfPrd
C3jUB25gjFqo5FRTdPm25rbvDksv/ODAQl0AYjddKkAC03ddPG87me7tiiAQSzyCRknjvMFhvRJI
/930vJbSgOpg+pZj3KCR6a/2K8ZTaqEmnvvw4Y+Dya/8umxbIEvcd59xax8CwHNaTyym/WOhAwlP
yCqtBkFgOwZLDShxKj4H2b1c0lM0AhC5LFtzuPRd5fZ1hsAFYlxN9DVSgT230GMQS7U3fXJ3LU6U
48CxGTZFjtIEbvhg4dBGx1LDuZtoZsuCrk7c+DG4szdQD0FfEO0BZ1nfqbCuYY3q8e7hFSqCq79o
Sm4Hl2xWm9tfXmgtaSaKBWTBX5iBZ4DyP8q7ksUNb9wwAoQXDi/FgUBIyh7K5l4qqwYKnr7rNkUF
CDXulE8Iing1vIJKQ/3OkODslkrZQ2+uq9TSdjwUqyy6/YSW06JSBKDaTkVMon9qm8jvQrVBPTKO
R3lJFCZhHL0xMuV8tDQnxvIGQvUMpBwhjCAJdd50vaoh+XT8JizmFBTtkp4yvlnBY1egIclyldmd
mKGbGMejt/CanmPmw7xiwDgopknUhBo4tYBbAKfNEmRxN8lZSidg1iJG2ljx97vcKyVK/6bb+/ya
Z0eGvJMDrnH4QTG88vA63UwvpnC+bF6cT6UaCjvaJyxzcfKgNQEAK6RN+gkVn7uvwcjyj1q6UYXr
F+8yRm5fKG5vRfikOBpkWh7zMPdwXzJ/wkdWHgiaC6HhkY/V65N7TLHFfXqzcuLG3nLUWQ7cSdpd
pHjSbLG/rYe9Uf41SL7MeiJzQXxckDvGpmA6mBMvBDQ9pVk2l0HuPvQFH1Da6x2+PYMdmSdpdYX/
96BGARHUNKwP9PhrxlnitUvIKSYoXXczGuQFDWXhqWp2dU+Rx0y6QA/DftNk0qWGIOurQjX32D/I
23rHCc/1qWoWYTLUe4atWYCg+vV4UrvRGU8SIqbEr5GAKK2YXf/8P+XUOKUGvoFo/f7Hko78TB8z
T+SEprUP9Rs7jj9rNB7HKkxQiKDSolVxGf6QhbP2JmJbX5qOldGJrrwhMzIv/UEdJzmWMu/mpSpk
c0db3qgNFljI3KElR5Rd4eyZwK5E9Ql/oVpQuLjLnh6Vso89yORLJauCyjlBN3zy/EgQtcPaHPKM
qadVe3k3UXlrUIKIozR/wISEWvMfW5nYzIIIL4J+O11e4tLtmLm6Oj1uaiBeCxOXF0bSZ04wbtJe
RravLIzKKT1cBaQ5yWvzvlBubb3BMYi2O5aZIRBTLhht8ISeNDQp+5BgmLxFfcDaFz7vtz9WqxGw
GsKVwbVAr9VQU6AwGBdF4gegYEsbl2Oh+xCxFOWU++Yo6U4STa2ErKvpd9/7Pc4u65+VwgD4qb9p
ox39TopPtC5BGCoQjZ1o5DijyUpPy+Y+xKc17xn6i2Zvr43HIYspKKmHlc8fKlsjgJkEmtYH1r+U
c+rNqgaCn0ZPv5Ccgz0p3M00Gu/moMi5frM57C+swmBl+FEUFxTu9zY/vUnTcD1yCUC+PSPeZuLR
0UPg9p3rQ2sjAs8QjaIuo9QKvGIbvuQCirht7mfvTjsnuUdY20BQcqbhzbpSTMJ68qXEehtTVObG
+EAt8bVIvBvomYPI+f9QIGVynX/i0pDT++09wWEoP3YDQuz8H0YFD6bb+Hb9APF8JnSsgRKnJcYt
Mt7ktPEu6Nwr4SDZMgeR/vU87L/uCFO/Xftr4K5EKmyLAnGH7GgJUMAh/rjMUu0Yo6IwYbdyMhb2
1S6hriRvN9OVbAQhBYplG6pu1BdQjBP9Qe5bmqgp8++J0OWbTJJDGtdcDfe9WfTOK5jpK/zP2+QO
k7T+mKhkK5z1kwHvWKLOllKARXH8JX6zhbaABQDioCr5ED11zmd+6s//y4UAKRFduuum+0q7Y9Ss
jeBbmRVy5URxzG8xOCOu5v4/U4DEyMhMSryYxWvIpY22hx9IJxWHwaVIxdLFvrHteNuOP3zckb9W
08i5Tf1iiajKxq8OQ3hiawCUNB6x6bXr//N3xGXUceBAgr4GV24g2c+viEEnHqPUOr/XTHUjtwTE
BPK9U6bbfH38CyVJ7AeCVBNpFiRiu5t+KqGQxQhX9kCkO2ZuEJOdGq9I/ZsmBXoLQ/oKUBU/pQ+Y
crtDovj9GQv4sd5Z/GrUTkCHXrs4L2v++It1AYGD/+UeGSva77aam1HZQDYRg0FCvFsSpga5DnSk
ur9+Xt1RtQS7zfES50Jp6Lb8hBxYyS1yzDAVAWReySc1c5Dl/N8sZ3WcYBT0CoXRlFdE64s83ZHE
vOdgoQiNKE1W08tUV53cc36GNCmIw3/gN9ifomTzPsITkdPY5fj3JarRiFBjXYDD6iTCzQkJ8RO0
Eq/IeDf5IK2oEAKf/PRcnUYxkeLeCQMB82w6g4pQ21uEocTuY+PWzrs1Str2r9c/nrASw+uXZMu5
0fL7qTXXnHrGagx0My1EM4281Zr+V6U77OQTZ7ca1aExSiR1DSr2WkHLus42gcYfWUVbCBkeZqgT
Nt+OP75NvhaCJV2k91wBrlbk/5BkX8AwUIddDhLNkYODkIFbM7hIoKtyPvO9K4vcQMUADtiPyAFL
Zy30Bf8/WLGf7+L4ydivXUx0TlDDWqTt0R2NW0Ab1hB80TxJIdboTefySt0ktOA2eJRLfW6Ridol
YVfExag+ZliLrAL4H/53U9rtoFuTrcPH3vqYlx4jITxnRaT6gVTaL80gzhHxzE0sT7lYEkcwrPIo
4jgIYoGbkNO1MdfdTvGzWzWLrBuzosOqtOcGBcqmt3/0GXweeoc1TiGTx7dJpzMvswocOpchvtrd
GLVBwixXjx951R1+1p/Pw2asalCYNR/J4SYYW+PW3dF/E/BxrFCmNf1Its2qHYj+xTnlGtL9K2Xv
JO6JrPAvaNVIH7jD6w22kFjYcEx6l+XXjiCkBS97wTKk/soy7BKQQWTNyvu1LR5gKYVZ7dAU0qIZ
3AeZdzRQq7nuAQyOYawhd6H9AgN9pUphKnjQ2C92wlqdk5dneomnwusDSyZxS9cwBJ3iH3yxG3v/
FfY1IE6pjh63Ko1hnjz3Bkp7JdjUv+CGOekENsfws6QksmeoG0Zcib1OjBMaUzpRniV0H0ZJPNpa
OSHl1tZL22tadhZIGR10tWC8NK4qYYq8H2V+Qb1+hNP9DkwasQ+R2tcA9qTeqbw4Syxmx8EvaGz3
JTBZ+cH6Th2KVusReUKuxbCurYvEqf54Tlz9LTZctOoGmv4Aa8ySJIMaDMYg6SIqGbK2NnIRCscl
q+nCqejxBYcWHPJLepgrRYfJMQ4LUxCfF/uR/Vn+BruISm0fc2KDDw4T1Jf0M4TOdp2ChMN4ZKWQ
EmZbefGr/yEDPdWO8EUdvDWfWMYSXuXUgtesPyhCjsB8UFWHyggLB1C1Arfwaxzk+NIsiK3Bd3jo
/dRlh8Hzl7ZRXwdUJiBcemeWf6NXi/724/+hFxSxExLftdtW4Gd8h1wk9R7k2hqRwhbJbsl4IPvn
jWuKtqGoHZqyrJxOOcYArzk1aCmP2AjzXxe89d8PIfKKbgkMM3H8jCMHx6JL8EwlBLoK+kd3/a+B
ZBKC9Eg7T+5ShhQ2FvWckya50BD0bAeC6GPAR0X8GTmmqPc5WkzDexs9cgyWk8eJc2ken/S/Jft7
pfz3t10h3oHr3dK0Jkiei2W+z1yKb6QyIa4xtJzt9lfqqMsGS8Igk6auEQKEEtt27uXfLsiTQlrZ
KEH2+Op6NKF+J+9thfBrEvtreRZ2jj19YKV0/b0Plx3/jBtxv3ZKsr16vwVCWmdaFb/GI9APwi3z
Bj+Vnc53BpnHMOGnmm1iShz0hu3Gh59u7c2P3JtXDISxyYbXRa0j7pnQGoKeJuI/zBP2RbgBN7Hl
j9vNQXJracj6R/26J8inhCpGuidjNeNqmuuKreXSD426SskUeTWbNaWiWeoAVbJtro5L2lSz5Yp/
SX6u9RdMuEZori8LAEJ47spDGNIkQsK1ng2+AuoUyg7pV2GOatM97otLU8zStoPcMo9Hk9XE1XZ7
odHzsS/iqtWYbvzBFMYbIJjru33sBk+1d/Yq+dmB3/bh1ptExrI1uCSlJoEkjYE9CviDJZ9rSoWA
MUIApvN5TD4h9XF1HzONExA9xmT0yAS/8yDcjYsiYs12UjCqP50P3LiALe469EiTBzNkOEJwLsIQ
T5CFEiHYPr7WpyyoZZdZOUJPAmWjzySgtRuf5JZFG63gw/FI47x4AluOcq4Yjxv6dhnjZh0LrGXj
vTVUMtVkqux+cE/rxmZc6phW0dQthWZVPq81nmxluvMMOGMkOtYCKIIm47tyfAesx1Va0TcDhfT2
jxTLgmXp+0gqvnWmg55QlTbp/dHbLtFL9vj7XpCpNtSA4Xz0bdqJtCPD6Ue3DVLFXBOphJydwQ60
MDaqHV8r/WNO/lLruWqW5Iw3LS73fHPwgKVKGfkGhKT5GAZjozC2qk27fHEcPQBy1phBUYX618pb
EovUyUlOFxqUXMEbFAWVEFUu+uMC6/pYYd6clLnDGgGeCOmwygC/vmZSedxYw0c/sGieDg3UqpSE
mciR6/hWOQ0Oku6ltmipFimUkjop+DxE0TSYJbXfXH+qdcWatzrRACz1pnD0qPNJZhuXXZcZeZdy
9XPuFGJThGpYSgbuAh9drnTsK1PH/M9ehvcH8RD6EeF+Ye1UE5ASe58XPsHRAOFRxogVDd7mWqlg
tCS/5iwzeFpJUqzIV7keaQOtQQwDpVjZCTJ64UmXocenmoMP/sufdbnEBeHg3xdHb7jRiuABWMRc
GBwB3fCu5j1CqbbzVnF1JwasHvLLSidE8jfGpAa75+VI0k5VdDV0LooJoJ9aY0L2MxegWcdlmCNb
4XzCqkvrWwzGsJCyWA1/+BySPNwabdVK6heDsEZpi0XeUUsvLwbi0MS+4CV6mtQKQf+KjpGDqQ63
ylGoQiioOAXt8dbjBA9+qdCxLMVugdkOokPQ6Sk9CV4t/Nr6JIMeDVEDzl8j9XTVSid2u6pycivw
dHL583knqmaZaL4bUhqSE/ULZQScdQpHT1RBuD5gdIWA0IqeWlbIdb5nzHLHQ230r1DWJSiV3PNh
1YdTCkaT83y3CvINxUT7Onysc05mP20nHz/NWGX3n9ZIhmi+tkuJq4FhK9zaEe94gbmUx3RTg2Uc
URObXidwgwFjS5qIsz2VYUVKODfDAeJiTlNBQrtEF12XfiL6KZczHOD7on/BEG9fDgET0IymnIEZ
5ewBJZRmH6A9FDoexxg7a+4WjxSyPS3hmK2fipd6CblKU4dJ9/ZNeHN+gGBINhMzAconFAt+DfgD
EVXq5nlFLFI1QXAF8LTpvIhsIe0LnbQgVv0qi1o5H2T/feVhn77FWLeL9KC1Yykv3ijJq+/Dll9J
cLsqg14ZPTeUodhqLRDWtrSMLNbdhB69St5KMNuQ80vU8BINODdiQUaKIL/P2sSHHY6Uecg9pUfg
sL++L3XrFU85poHqC6TlPhstE71ywPbkSbURCMqveMTp8eKDHu7KFrG1MgaZc+K8jef1Ptb7sn4a
Q8bIdW3XbWbPAndssF/MzlavtDyuucpmia94u3eubhi+laQpa+7Bh/+5lLPuYBLCQce/z+LWUMm5
eL7Bzq9Xw8pmZp8P78T1FxXf1rKZtPcIdUUD+dW5vDbQcb5M71fzn7rGEKJN+sprxg1UKlindBLH
XzZ/HDXWb+cVw5rJlDTIhRWeJez93BGy8Gkvf/i9ux2PUImLYDJoqhrUjUruh2kctTg475ntwSC+
gjiGjZvRkCAZT6Ia7Y/OV9HaDfSD25i7XZ4GCmvwOGe2VR1wwNW4wfVSQSHggRT69QdNFbe4/svP
jGlVlni0UaWwIBdr0C1Zx8DQTkPGfwtonmuZXStp2qG1lW/WNmMLWaoHMUe2VAa0dRA/oMaq6Ji3
c5bN9Vaf59WupZb4o9FuAjDxH4QezWHmTTu6QuN+etUgXh08J2QiOPEP33zvMlqK2gy19rccSbWS
htVKvtjguyr2EXpj39YrgqzoplUF6kacqPCW4ZZREXKD5ifRGMya930a1nB22TpW9/GFjPm3oxUR
0Wh6L9jz68fd8baFCredN/r3/ynASEo8BW6j4S9Yz6LGPbETOnlnxklTQdGqZp8cCQMP3LykIc6j
eJxnPsxsyPvpGWUHFHS9Mm1kh/Ki2K6oFmn/HOgj7RGIZYjL5Tj1BWe0xrJa1/08LYZpaMjic740
Thevdd0BwapWycHNnOK/wGZTuUlF+9L4we/LJt7HfZlcLu7iaKCtFMil2Hkl+KToeNyHNj4ERY3E
Y1x2PDN5ublPVqUhCZXmZ7/bmnFaFDLl2jWFM7UzMN6ND9FEiYiI5EHtNVRn437z9icfUMd7ZIfR
Kizy7eEC68lGKxTr0EwRfH6oJFrHtAW0viAxKt/McMqW3maA4Q/P90f/SdcaOyfw6PqxDTbnpY60
AZet1faDbozR0TS3nnmsn4aHD7zhGRmlWRwZ9FqxCqpsy7HQFVjurAUCYKI9ukKCGqmijhOolowM
RPH4JNUtxN0ycPPQgDXGn7IXPhyHiP4KVCyL8ZF1E852EVUH2wAwJriALXI44YHTJZX2TbSdEdpi
8ZosQDN+0ZFeNitlhKlGtRb/rCLnc9n8+qokeSGE7B9LDkosbY1pKHB/jUSajXgZljTRIAT7sz4F
s+4V6cA2WQZWovqqBCdIOc2TABUm5We54LkmZfwcyzpSX9dIdQvTgokvKHYCaXUtuD18omQHRHeQ
KwiDDrAittZDlfwqRhU2MvEZbdlElMAhI2Wi/dUoPz1v3PHNhjm4vhxTa1w07oAAeMTeovCRSp5B
0F8ut5Jk3/EIVNq7S1d9q1cmd0/EqLuD9uPKicEXzOpy2LuXpxnDiWvFPw2Iy7w/8JQowYQcMwJd
QVP9AovHFQcNtta4Cd9pjmCNu/31ek07KCsbOEMoQ+YF6y8CPRJ8lXGtiG4T3bNqLDjm7QqGARFy
jO1ojUsd7kSPS9hYILB4cXfI2omcXwcd4/o67+OpkiMFj4eoAqdTwb1Cf2K7zjQLL3FcCdc5pcbJ
/MVUd4qkEMRnN+xVidvSEyRtUcmYlVjJB7EDAbVVq+tggKfNJjuTf7/vh9VdwaZjO9bfcS1KL4UH
h3zPl6Ifo7cupB/BLBiP7mxpoNZwAf4SL14xFPMWpEJeSVji2chRo5nvgu1VNvBpCUwftqizcZ/m
c1movSAWgCn1LFNzj9VNSYnaUc3qzztHvfC0MuS3DxKaCFogRsJELhtrx0cmE0K2HS9N41g/F43t
WW7K2fxR0oqjfcjACoRu4GhmhyrAryW7VGINMyZSqt8nwQpqMTXgNzE0ez043hqBt2DTPykxtL8E
Wg7w5wC5HfFU6UG/MBbSX1nJAvotr00eYqyi7lxtbfHrd4JfwGUJ3Vl4x7D1tWfSR6ZoBaQuYlEC
PpRe1vy7UZC/xz2s5sx1nYg1HZhKpp/eQnuj0XKyl9icr336k1A7X5ut7LUz8A4gKzgYDISUiIvZ
9kA5M4ZJEQoH7G1nnOGc/BteZemVaMqCw8gI3L21sM7dc9cH2zGH6mfipYy+PjU7R37l02oujP4Z
xpG/32J0gfc1nLPgX7A6NfUU1DhA4cZpYmH+p/Xa68UbjF9Ot1aCct3d+sf29ugB2H6QrUnlJ3I2
jAeSEzJpx/e024fQ3Zgxhg5WYzbaRAGQ8lqtp95un2mNgx4g+3oGmUFi3++eszNTTB2WXnXUz18N
pKOI+SQAEie/YsUJjIOA0Oa6zDaSgzplo0kFPtRTexh+luKacjw+JFgDwm59caVf7l+ZZK0FMHBx
RimYgqi24cPZJmG6aMGsJlp6t0Mvas5iOhne1JPbz50rfR6AprSoiBAwA3xYeZBqKqxhRfMJ8aed
iLMYFcS5M6DI/esUa/7tbc+ekpidrAQ5QmtuK8GJA93dIM8W3Vihoqe+wZfYn2taCHIOahQ1KOoJ
iCGgnJ7H97eSJT7gojT66Bo6uDSUZpXjGEs5Ve8MwyhLzwMqDfs+fiCGCwycdMHt9D+7OEdMA8Sz
Rw+LnbZ9be9aJr21K+2pVg0F9I/MVAI9YON2TVvGDwTd769s0zJDMHahAweQGyv0jTbeFsZjjGdO
dCJCu1WS/TZu4vEnkCrFgHqq4V8afcg5oUf21+Gu8X1Q7+ETLntVMhX3ceFjmB3JzAiAM70/MQNG
95fZaleuuRxc5wR3OdUJlOcio+t/2pw9C/6gn8X4UL+W2FX3fl50+04h1DE79VTGdiiS8yFaMN2E
fUrJ2PRrI/JDFEyaSpQjPeshYVNqjVCggPfvm+t45CjsW6pIKOtG1mRAFaP1Wy1he/ThH7rJ8+Th
IR3lQMAQ2FTVQrmKbwzg+NVFElLYmdmaDkqJDFCob7q8kVpiZ6fd/0NTgr7i3S15YK1oyjdG7hN9
74DNlzOzX2+myBxTcZ0sTT0TxpyncETuPm7vxi2VQ72cWtsjcIelVSraWJJOj8Z4LQUz3GLuuANj
C3/7fy0ZwVcj17zOTyOqzsFW+Jj/JqKNOxsPe3Dkb4D+lM+huQ5efay96iScqTpoO7jbp5cXzKNg
TDjW/oav4eF/HjSQb1449WvgN9rUhieUYeMFeUyJO9VgZZDPOOl2FubG6hfKCmh2MRHOkGfU8u/x
ZPG/rIGMXpYEe9Yx9ylFttSe/PX5f+r/t6B5UlwNItn2LNiS18QKQU/k4tLh63bXHTpUOwPS3YVL
z7m0aehWDYKfYLS/NlI/D8zAfbbyurHUVUzRexj+/YKCNkQHnBVNfmxurE2HdfXBDL/rQBZni/ZA
6eKnq2MlTRWR1+Y/Jv1MVOJZqqf+aeaLrzFvqZdMxxstqnuRRekYL8b1q7qHurlYp9YKO4ibzSmN
qZgbytnG+emaRRqYMRRJZCackG/e65eAAoEz0sWeMpDI3YAwNLs7axItkckeIbMHG7gvzhLm8e2r
0GfDxlDXwIwFdlH1kmEzCjsPr02Iyfteorm6Go9pAiM3A7I1XLJEkB39cRb89Hrr6iaXzglX7rTg
mY4mYaEvI3EvjQGqOPFBRr2HXbkSORbq6EVE4ie4bkhVl0RXVxzfnYTgj+0P+oXgJN3Si7EIEZS7
W1OlYhTcEoeO4yOXzOOj3/HFRVRqzDLEySSenEQew60yzEshB3GpcO+2cj/ffPE8L4gGg+WdWS+p
lJ0pinzafeopM4hYmRIMMMaeE3ogs5rpdxQFjF8IYwCe0l7sDv4K1yYwoix2MiCnMD2mWA2T0+1C
J3spQi1iUyZ592jQohMzgvTYGBW5dI+ou6Kan5hSnLfEzEuTyOzw2GZ3FcNK2J/fREAGi571cG7q
rWGlzYCclYe5lAgACxlt7QTVVZZef3Ro16WioK2nsxpbHfG2iybKsewg9Pu16bqMyCojtV5AS4sZ
Tslmg9GVaWGRHSbFRaDUeKoPdmgv/E//j3JDu0ulbvh1mcd2Lag8pff0IdlPW13+Ocu/guyTVtAG
M4vRFwQFc8SfVUur1k7rGRV7ur7mX/5bAGE7Otpw1XV7Wldgq9EpHfshVAHbm8KyrRr28/VSCzT8
z/5EmzWPtYfVzQ8nbPtnqTGDxQg4D0fv9jzTLNhcK6gtG6YEW2u/i0EuBAHg67P6ENZr+fnG4mWy
rHhLoJNiK2eBz7buF67kAHCaMc0Qk65XCK3qIQ+Jn6p6aJde4g7Kc3pMDkr+2dB2e7NMIP+1AB5L
0ZnhSbAFLQOnH4kXVcVaZQoR168uws4SrN8WL44JfzyJcpwwjXSyIeeivGqPGHVX+texxCSOdYRO
+CTFyhP4gF1E/jv6++c/IUCnPZvcR8ckgCAum1SMt1mWKWDNMyRyQHGpyDKoONYTum42fKL0fb+8
GlPdNKVjRm0uATOPI6LflKYH01UmdqvFGdiVSxzN+sIhXOY1rIkVHj4+QZwN2r+z1vcQ4IOS9ZDg
Sk+tt29GafArWet2XE93/U8DZSkbkZeN2NWO6Dt49BQWS2IBc0ua3yNLCrbAsg1bD0wRXk0e5AaZ
VyCTVETurvcN+dF/jGeB9iKNUri5cTp2A2x7uqAylXDARFiPvVuAEFECvGFRHfJ/tCKZ/PgRJ6al
F8ny3A5HFzwJ17RRCIDo7hK7FGcucFrA46oEy5iG1nujqM2SD7Hdo1WfKm94MSRVda/yTTJinoe5
Ibd/w4Vz1Z4TvinI5tV2Yok1wIQo/AR3n3fjAr0pHiTL4XFkXM17F6yoHURZEMlP1+JOPKCy3fcs
E9i++EkINSG4CBtvEJ74h3ahaWF2lZwKcB1skhp9DdhYHcY1vyx9vsyQX1Uu/XgkR7WuO+WrMSk3
nl9guyoIDUGTDRrjOgo4UV3Xmp8QsCsok3PScpEo661w/LItc8b//bgBH0zrooau2flEQ1usJgAd
zuhxqyplQ6FKFmgRow2N3HFB0UYzcUpzQzDXjqxF8tUm3lUhvZSpET8VNV440On17miCpKgH26ZN
p52DGj/huPvn7LpUkioYDgueTvlMeX81bG6EAA9JGKouwy0dwtcUIhsVZJQ8HjKHt0IQaDPmbS5F
vKYpHAMD8HJ6Op7fvRwj/XYO2nV7mBgibprwSfRxBXK5oGISUG75cOdVzo2meG5x8k1Jp/PZT6r0
bUYuTkOzdiA4cxbBTzoCWl7TI//Elv1q6Swdu1dk2bipgRp1v7RvRYR9LXItLkc0vxZ+EQSvVz31
qWuTUc4X/z0ygqKjyC2CAqpy0UJcfs6wZZfE9bh9/6dOyQ0TBTlxEDNNPGsQbShGq0liX1LMuZZw
Gf7sVPyxPcIWU8ggyEkYCP0SUGOzJgz+UCdjlacpEyu1pdu5/bq84u1Es/vMIXd0mcmNEga9XhFK
rEysgQmcrz8wt5n260ngwCw9WoJNDETsVtdhgRRDPgZFkt0mvux8uj9ainRbJwl/Q0bQsrghq/mE
3yaQpGak9hmBQcy13kPsRWX1RW1u1xYuxsxud4oXlyPZOKJpQXLT6kITdLHKDmjXTpAYDtLBxlc9
pVoF0VGRn9ghJxYzxdA8ypowWINSa3fWPlYfOzaPiPBfGApYQmdbqVRdvH+DxPt0lmMWJ95XgAo4
w8gkvneTKpPLmU8IW9OGEEGF/yPo8UO5cpScJSLyDZd9uIF4p/sUUeZsAq8kWxnLjjsGQWRaKgZj
telbMSIkZSfa6Ijq7c5WovuHNOZyUNhrc6eEd8APfdoSP5bgDSD3kCHah9/nRl/tL2DlZtug5jEo
+i0unrqSEZHaCxUTxprFpww01wCXZ+eUQv6DTTIK+3pdhPy7LpZyeQ1vOMswWonOU07ZXoTXM+pR
P1wLQD3HlmRrHuG7dO3iUkwaIXQjxXV6HeZt/2W5hRWNTQwJ4hZ4Ej8nDZf8VMAErpHY8HTCtw6Q
fl/k+ckaiCDrHbCoBQwTfNO60OwnE0V5Wz+oUsgur7hraUxVWV9h6rtRjW/2BDVoQfogaocGHcel
YCSBBavFRnHwls/IPiD4uwoMnLOgjSgZhoK2T7ZQ6vOAcPZezeMwwDY3ipnh+QtMcfe7qGrV2eoJ
BuA+AjK8Sghog1LETeNipb473ZGEBHDr4dRqW1eT6SxBCpUFV9HWpbUGgIzpPwlfRBiQoYMcA6SV
KzDHPddBpDW7/+iQMo1CkGJ/JRO0upsZGhuYORjWAUe7UsAbJT/C4Ib9yMZPm7sF8D4kZtiMuy9X
NR8O4IZRsef0nW5LYAHShdt4DyDu6hpzx+W03zNz4Tfakhp6h2x/CeD6Z73cRFTyesK2kDu+O2kQ
1AFsUm2HzRw2ZKGajOeysyLrgHDxMCzCZIwnXCSCm2QVL9J39dtixNQUXpW1uXDMMYtNkT3FqNoO
Zlh9bajVfYOmKZto08/O/k36uoJa05Q+I06alvLkxsb3iQQb6iPerHesOn8xgFytOeJdQ0qpCs0T
yfFQGSyqZV/QukVlSkF+nzHwCJanr/0vJXpq7610iymyjq1IaV/NYdThVCeM6mf8mG94HVI44A9G
Qen1McMR+I7TK1BLugokKx3+CxNZsXtjahbQ06q0uTti8+de5wrLQyjhscmNHC9R6fddc6jwWvOM
19KqMWqT0NlAXqpnv6w4fixLuBvxft3U7oFg2d7+DtJ9BbvalHuh6dNZzW+H8wP4UVryS8qKpMUE
WPhQPYE8z/8+whgSbh09wlZjQok0zq/fis2QZQwf+ybMtlkr8kmUNe/aOwZGAamE1GUUbIV2F5AO
jWgYxaYHJZfmbAFGdj8ZshgnNEaZVuelmWuKssRybQRckVtgIWCr6DMH938BuvsLRZFp0Pf66Kpf
fBt35GUPz/W3QBumg9a2GS8GoPEj61xU9I4fPI+/R0sOyAyFjZFMTzqoKXDD+euorLf+QUJLN2lY
jfMSxeSsEjCdCrrqRzZTk0cnx7COQAl1O0aySeegY64/2IOPNZGk/8ouJQKNLcNIRwv2VyY8nyce
uxlAxnUQ2j4K5qa12291R7Yrrzl8bUmUrOFYw/5QjpWgU7l1P6wYxu12C95ss5b0rQy/ojKnQwJg
Oyq4y25gPpiArAVYShCJ5MXRGs5hYec3dCtPvdviEM2S0F+TOWpIQpnDSxZ2YleXnCVtlCiJjF3d
yIO7R+ZNsMpfDwhXf7tWfOkKKD7W+wEtN/wiiD6ohm2rvbcHJJcA6CT/PCPLfRwgOROz3+y9jRsQ
ZG8DqgKoU4s2HRHdv976XISGW8xMD6z553aHQaXp5xMBS5jXUJmOlQi+90YPUdxBbmGpup1luLfU
wHgcov0KgGKbq98CumW8QSN1yi8PJTv2MA+8W6OCuefaL2967N4g12J1k8/qfc92NusoqcsoYJEZ
oD6WqoRIu5fL0IKRkauGWXzSdxH5+UthnGlKuNFqdms3quuqYNHd+hc6KTx0xTJwNk8INuV2NT7i
iDLPe1jMn7+9NSW5Te5VhhwyC/5Nfq5Kw9a7zAcVeho8KLndyLLAhw24dUCO4h3OA2afB5liKzCp
XYtd/Wv0T2zVe5xIw1ZRR/zr5JNsdIv3uyNtXTCCTCdCsgnvIs2Yu0i7YQAZanpGONqGdsMKDavN
yj2kJBnv/wnVr0jK/AN1DINPdN0Fj3pP/T5Ka1e975g3MzOcktq8ioONkYgG/DC1Id6ASXX+GEIH
RgZwgI/BcDwWw3DgCU8zX9bwMr1mfg6jv2d3QVAxI2c9llBsDEEnXsWOMX+VMhIBkeM4muzd6kZC
DM3Eg3mOubzT3PLFbCrsedy3Wg7zf4aO9sFIDVuJ8K+Fyk+iCDF1REqmSLVSmGPwKPIbI45g7tTm
0clWuGzbxAWOFBUB/jkwnp+E/BJwBn0Td+rzkcNgIXtm+w2WJ+AgOkuhuuzk321UKS0zFslfF50Q
iFfEdRjfQv1Sp0pdN0Ea9QcY5ACVLeDoAPcvhgfesjUOYAyaA11hEsd63cmRYyHaJINeVfSDdEnJ
iwJ/ILJ3GeWxHdx17yzklshQ/3RFu+EP/TmvA4BTBwy943Lg6YCuK7ejvgve62cJ73T4cAxafxBo
wcix+LIOLO2WVfNTdtha2MsL/B4545U1ozRrto2aKIPvJhcjLjxpLNi0c6jkS7hZGE1rTq9z/Dg5
JnhJL5/sUsSQUAIOEGk2TESVHjVjbekYRqFwmTlPWpAogat0Qtyj2xGG1Dk1WUN/2EbsJAJezjKQ
3sAX/t8RzxYx8oU2ULMdATOzjc5ESnuDTPXzRC2i8JToJn9MQum1ree9p0ymxamXuZOx1VxbNt1w
o7HzEgSYcWbtuo4o1GFYT9qM1ZVDHoU6/PNuzNaWeAW6K17v6yW/0sXXIedEyxOV8VSidkR4TJFu
BwfHrfVMF5ARNMXPi7rL/A79MWwWkTCz4KGv2qTycRJ3fQ9xZLzczFbVZHBc0lBq34AiyofbX3ps
8vVjCJvySHkKpbuRVa6dVlIt6W0gnPgIe9tOLlDeCd7CVnjUwYzzvaQoIaF/1gCX4GZmdiJr4wzS
3SlzFOwcsUTDtJvM3i7qa51agdpt/CP/we1I+aA0rfb3UGq6O+NXupajZuMYj2R/ORXib5CORW/A
iUr8X+snwoWOe3RCxf7lfNUiymEWb2yP6dPY7OKHOVXUpEzbxJuLIMGPGlYQZEQjy5876+uzp2od
spNenbjmlpeFjOItuBxHLAY1rr/OsaMpXHp4u8uMhwBnmW9O1qh1cHPn35WFhAuCU6n+8ms4HKGh
mkZAntmgV4SXyK1ONs2k7g+5M8fUyLScutjUumVDG96NmVBZH/TAguwOXMcDsykY/4cUKpSFJHEd
XCpvYo2aVSQE4xSjDUZ9ZnnioT9chPRJBMvRTeM00nKEXOxfNam+eFIdaAynA39yCZyk07hTFTqM
WgErnTK8VT8bvzPasUpcuI9fmNCpNP+J1vo62i+olvoXTx62ENrk8IMUweiDuU3821jdwqpVmzE8
4eFQF/CTItISADFWjz3nYZqynm7MQml9xKU+6MeZ+Z1Mmb5TYN9fW3L6yTxttXmErMFk6iTA0Qy6
Ae62IVVUNbRlJtA97eomtHTCIYc/tq+EkY42C6lG3qGvqK7SOzky3wOu60wzc6nRYukeDc6xUmNh
Hw/Hs9T8x0Eb+H46DNra8TeojBB/eLSLLcnJht9++fGcDP8H9mzGqwYAW0iXpV+8UT6vBWUQ+mIv
3dzU2rql0zf+6NqMmgJ0uI9A3cbJlC4ORcbecCFKHICbOwIPzmCjJEXV3aAxyW+ye/hTt0YxQs7x
3RXoQV2GjP7W6+7EMUBnqn7P7oceXy1HUOuvotk4YEw4ebcOHu3Es888EqqXT3k/no3gZaEZjeuk
9VD6GWyofxtSAAp2OHVw3IO8yBPfaJixwo7NqlqZ+LalwmiiODvR+/G2KizF67/VMreO6ZaZd0Rn
Uat3rA2P63Z6ORiLgX4V5G1gjGuN+8jnqvaYOU7CmDYthuBZ5/7d5Wc29xK7HcV0WXJteT8tv3A+
Id52oPI4mLx86A/UBfYiEp91f9G85sJJGmCJRRk3L4pxnDmshndb/aFyIIy5ARTZscJbui5Fx+vU
Xyo0wn+8/qbf5KIf0cNRIm41hfmhGHsEerztvUXYPXWl17nZM98nzOSBEzk81WuHULoV/kNCGm1W
wv/HPAL1TIHloip2n49YJNJGMDV7C5GDhO/axoP3sTq2hOkYIoKyX0fPeYBW9r5bHoIPnjW791Qp
4P2urXGWvewqyPYHbu6Zz2YcBlH9KJS65jB6I9BOlKGXREp+J0EdOLfUBQnne8COdUro7O9zu+U4
d472AU9aw9JyJCJIfkSt/uRy2a3cVxSfVy4du9k9BC8PtisFtVh+0hyH4DIS5QoCEDvvVg/Rs7KZ
SeDijplVXPXmqeH1Lup9vlce/9tyWM0XdBhGPjB9vi3EGwQPKKVveMoBF7tn9UqAKgrh/CJdSBR7
cuOnSt+RdzflZgsTQU3jqQGrTGwVyMAbbcb0qDJ2beF7kuxKck2VFceoSzsnCSFBM4ImkD36OFoa
Plj2qb5t7hnxr7B1BZ4wwSUI0FK1JYHSxkknoljLLpJ4q7zjRBZc1rLV7bdNKOCzjAwFsErv8GZA
oxGsdLaMlxLxIlz3BONCJ0eeRMev+Zo8BZjhKWLEz8ZzF98Z84FR28NJHWERiBBIsMJYLUHztrzF
5TofhetbQ+En0LqvHl1yAQn/85LXzl+zboP0P5jFRzgxoMDpNiqQUmu33ChNq1kACsOkJ7lJ1iqa
vTVojgN6nT3rL3fRfWU4EMAoxcUNiN3VIJi9oZ8++966iAVoXXWpKH2ustyHe5ZqxfK4zdg+V8zo
423OUAangbDReRft7Bfri9oevxhi6ifAjLhE70zorCYoCgCGMzoxJl5ehcpbYMfs8y61Q427I9fv
LxRL3m/ERs2OTk4MMulu2hni3JSP0GNh8tqO4G0svQm2u0UYXUBr4G7te7WBir2SpBXDUCDmlf72
uvJzaCeXcd8qkhJ/KU+pKsuTZfzAwq3HJT8hPYrho6EqLLSiDLQV3bkLz/B9rpYySfxSPV4giuaa
3QRZq4mODsu5X1PGMF6ZHpMSIexBHOeOSV1Gg4mJjaXTg3dPPH6XfyjzdoLXXBDrX5AOlgRFxr1H
KD3TElHXC7rjO1XHsKLJHgIwBARM3BTuMQMgsDonSpRG4gY/ru7pyuv2lMWtHVU32pELt4qnZiPg
/c261yvOhL9aVb7A5XCgxcZMtvkqrJRg5X82OH67NB94FX3Qnr+MArlE11uTsGFv2eVtwh/5BUU2
REbFnt/eKuT0XxsnZJ7IsQmeVEoW5r4vOsShyFKrYVY1ELtx6lkkl223DxAeQQ9V/ztLdYMrOVzp
G4h1f1d1ScVs7cmoo2lJFDjz05m+CcCMTigYK6CCUVokzaa6IldKufFVpuEQnZXw7DPyNAUNlEGw
HenaA7DDNYSVBcpucsD9aMxMgm03qs+iFtpV+FToGEb6aSyORe3HVZdzF6+UEjuqjGlH1FSoJONU
51bVGffdLXGXoxHiPw3nMz85cdPeFq+dDxmTwVlHHu1VVqu0EApMTbJRdNGNNuselxkeB6FphnzY
J3PNdoOyWejGxmem1XnfBLPtRoY1+Xs0t7/MfDM/WiZSNSqA/cdE1u6kwXovdifg3btSbDXCGAgs
ZBxf27XXH7wlyOtjZxO9wY+Zh7UNx05EO9Z5YOiSgrbSrUudn7g32pUe6JzT+V9wR/a+r0m64RgO
SOxIiRwr1mXJyLdBriCHz45Xyfxv4RmV85jYQDrPNzoZcmR1Vp7WXS0Xpk0q+aUlAkKB4YVE2PSy
/g+l/JKE1GOTlLJGttSPkx8GtFexHW35rFNd25zBurhYe3cF1eG7QKIEIYe0cQesNt0RlbRIwdVg
DmADEJ2YVxEm9A01Dr3BnRzrKqZikNoyoM44ceOpchlFgfkVCiNdiHVEL7rejfFrB6pk8v2M0igN
uKvkFmNGiwf0BAO7+HDYaq83f7n55GoZlt4vHX3RwyFLLPcS6YQoCpEaLq+wgdDKJC2S9obbLBiM
RbQN7yIhsoueXJX+DGlOlIWmhWGEMwT2BYFX+spKjwZMHpTndPCikHBkNf3e0Xf7yXiQiykqDNbH
LU+DbGGxfL/sTiP7mSlrEjLY5grmrrekb2yW7vFAOIaRq7IfdUSfbG9GIKmZEQFTDhO5p/ljyvgl
+mBjQEBNr8twShkwb+CxKnoZENgLJQ4DZMBp+lFK5zpMM0W6BOmHGF0/mMvxZ1dxsC/4IVzNPaCD
cYN2SXnC40yCZC1e+uu2LsZX9L2koQWTGFf899ughI21bGO4DJyweOp7apvn72rlUwAbarezUz33
owz7jQY991p24jJDAFnnQRF/hn1M0Kyg3Jkykrwi2UbmCMfrPyzVbkF3rQQD+fc7n2qsLRjapkCQ
yTcsbpa3KHf1nQN5SRHTpokYGI7rSAtLrlh3LptR2nYKOZOGimGlulMWvLClQbNGmVN7mIpkRf1I
0ty15hyUze0jInTrLdM743gaZ5oNtfmy0qOwsY7DCYbqRxayYXwKtCS3dK89TNZQ4m2oThl6FXTY
cZC6vv7lXVpB/hOPEVy6ijM0z309skvO8+lwn7AzOJQruOPIBxM8QfEua4cd5hHH34mT37AT6dMG
mAef4c6F5pJPc/UZGcIzuqsrF1ouP72IiOeEMuSkyme8XE+h5rY42FSIpdFQUqf1fFTHiL0A8hre
niHkxkbLPU0VyIcsBAHZzhzPWoETPwaFrDAY5QVTOnFJ/vKIhgZuM1TQcuw/83XOfFwhOMCqrk1O
XvqARyyZxlAgtfqk0FKoVhQBa0SMHl4x37l+dyOljBHmgSeKpH06fOL8ZL8qOIshzIg69lEpoLoc
fgB7pcuHv9C8PXyXtbnn/+kwP/wu59gEojB1PzpS2VLLWYQWWl5hYx2LvJf+s0OAyqhdS16ycd7L
+BIOCoZmxQxfob2pWODYKEpRubY0+VrQgvf8Y36vmx2T1UCb8yaeUJ5TstF+uffp8jnewS/RjndK
VWjeB2/ghzclgi1uYZmo9QcW0fqzZiiQbjIdWz1IgQxcRZvGDRm6Q1II22d83QlDjJqXwul+66N9
qt3VWD4Jqn8Wd9b5RJFeq9mL0WdHnherVZyoRyiEDk/i2s9r0JExSTcp567f2LueflK/JH87GdU8
vXpbjNZYsE4V3BefbglcCNTBD9BYwGl3ohjevPv0EumqpRpHHThJiL4m/VbaYSxdm1KN8xX7Iyds
IRPiKr2VZGbyZYwa+rY6Z24uHj/aSCzppsPnhpNHAJRI3KO30+y7Kjn09oVKCHNu51m8nsBDhjQ+
GCu7ZfSvcVy8lxM1hyYutVd0N51/caFmpOYT3NsfSwQfQQEtMj4wEdUqOLHKnx9Tm3jXVTIf5dWA
pb4Sy0KSA09IcgsrbwxM8j/rhJH7Ny0lq0C/D81zH5py7sDoVAvl4OdOwyFUeNA8cwyot4QvuUIr
8a41Af0Sj2OdisVaa+vgRXynPqUqAB6DzjEC7Ynl3osjB/5iXnqDGfa15SSEwpyPszzm8yazf/Pi
aVAP2QqRFI8pT/td9DL8u1PNopXi98j012krrtCWVjbLP2IEF+QYC84/HK4akROqHqwvALvZvis5
FST9a7R1oJVYPQJ+D+Du6tXP4GdGQyLpYdm9oecfd13NXxUsQkowYeQd/Bl+5tPWGp9EALb8T9qU
Mwu2CKb8N1BRy1fZkC8jtwvPvM78K7qJ/njHugCazgFLGz3pH+vQSW6C+RnSlG9o8rPEMifrdTfc
EPtlThhWrO9zuoULqnieuW0xMooJ9Bb3bDpk00hkjOmeTZw7VaWFjBPxuPmxPnoPn+B2geib9mJh
BlCwCPPtwDPazj7FLaC0ScKgLIxyhtu+GQjr4/uJSOGHobTLDmH9muxXT+A20j9QP9xJWHgTYBWd
qsT8HBEj2jJFcHwxBmxlv9CxdCD2PT7yUT6eFvquTf/AmzH/CIEOlrOLfazaGiEzGcZzeJjqwKVN
DJeFqwoXSNPSwCHV0rgC6zphiRUChr0CTLXKGPW8KVexJ8M2q9qXPSYDj5RIBE/V7LrRcYmgFKbc
1jDe5eLo16Wk7fi3IUvD7SBKcDeLHd4ocUgX7ksuWcWqf2ecrZrHtSoVa/uJAMAidbMx69nIgmDy
CpbQfvLfFESjf2zNocxl/u5yskjYtDLlHiROQtKMOkWGZYPdkmJIdzG+f3MPbLGF2hZZlSvofYxe
Nkw6b/xwqCGaakGccshKZygct4t53IBZacv+SCHxLpnAwmGsXJ7wlC/7Oy2SCXqEatfoywBfyLm/
cEGTK0cybw5O8hFrCIaAnXfNegbYnVkk3Z9kbs5y0HOlY8lhAnuu8c1aekmWpW2lAi+J2qrAamg+
UHHKUqHui45P4/Z1zSOGu+HPGeWhQDWbgQOs2658t5YxaL/h86uKemK502L4kjgLPm2gRUX8nBdl
3s9WfE67IgqDqGcs7QvJM/neH7LuLr54RdNJoky5Vbn4AcBSEuq/gyh+nWKpTf4w/3ZTMDWAze1F
Qu9NvQycDFVuZT1wqMg9I60y2sf1LAc1bgJ1tMwZ+7UTlai30KR5sHN7RtnGBI730l2Hj6GGsY1/
9B3+MeXPvqKCIU0Wtb7vuDm7DvY1ONF6n7i4YNTj+7ubm/MmtHADz3eMbJ0reIBk2p4fkusRReyr
cfNEe11huIwrebIoGBFaLN7zCR+AVYt1+w4bEYr/GkK4cNJX990e0hoTuhKtqrWmJRWnNfPrvyvF
xRl/FSBg0Agu+vndvolHOeDGenLA86a54LPF00mheFPbTJnshBoBhJsJ2CTWPqyehvi5OSpXenAD
N+jg5y3lOE9d1Rjfq0YR96N9rfrjg+mDx4kAaSL2nZc4mDlBJVi5VSjSowiUFSj3B7qHNHl7qIfh
LLLAL0pJHThWVgR1t9fabCmlsSNeu9IdECZ4TpWJoJeAMWO4Plps4E1uI3e5tg+JQVQE3PlpI5XR
hu0nIWVFeSz/X47PMK5Xk9ENqg6GfdrQv9Uz7dbb4MGMEVGHq+iI5OaVNrHG8bV9JFzb3Uo9cNAT
kLRSOnYf9qUQD0iC0QWC91OoZXMCqFiBKFynKV80zsHWKXRPNBMCZDhzDiCSc1JGBo0ksH1lMh1r
sn0nz+GV1LazPFzHM6qVUULhysq0+2FgHT1r8TlsgmG/0lW+Fsj3t4IXRScBvISXofxbhRuwVh0L
Ql5kWUzeNF8PJEXaeNSgM75yBLLXkf3AEfV5m9lQ4EvkusadRMrQL/TH/mUgIiXiWsTP8L329V+2
HpBFNiet0oLcEgrU26w2AIYDQ1hBxhqm2yJxSV3lQsApZu65EjHhavjJSLSVde5wb2A/pImcF7Kp
HLmVLZXTgEysN0KcU60jmWfgj68V1+3DXWOX9D8+UOo2xbFj8zBeE8ViI1W9/o+T+kLXK/deHXUV
dngF7L9D7+kw0wVpH4blch2ufrC1ltdb4XbhDdMyyO+pe+D6gz010Z6BGVfnT9pqjpkNNLXsaSho
Igxee7eWfgXWg4X5tfJtN0A4/8Vn0SzFoqJOOgcbSG4jxAjRnbDvQIYsMedvF/t4c6KZ3g3D/rEN
AqIuFT9LKhdzL1pBSNRhpQGhDnI9P9/IKP8posIrQDxfDUaUEJWbHqMPGi/BMROIbmcW60VnkNGg
aIhPaaGAJ/tCTywXvxn6SlhhtrgYoiSkr/QIe9f1fHvSRZ45G+T/cWvr6d/6yOxx6ytS+5vVKUyw
9fZ3fZxkXRUT1JG7o89uPaREO/cAvYBcsrKaP+jX9sR2T5zutSIvOp8lFh3YSDJ3cnucZBNKx+Ko
q7eDOq7kPZGl4vGdAlu8UeTQ9VSOkZcymFrBzGdS2o5BX9yMSmCOR6Bdm6XCwRuPTSgqJDMeDQKA
iM12o+R+u92ulneQUN68HyGVP6CGhU5JZyDOe4nY7ZZQffYeynmrvsCqq2jWOfOMhktTK0iakIz3
PGCcNnRRrr/0vgBv1x/meTAAy/xlwyvqVeK48A0D4uDL6zF1JcuCKtU2Hc+4H4v1DHP+UOL5k/cG
z553/TeIEo9MhoH+AZpPHz5rqyYn2Z1hhNTjREgIG58jqU/gNLG65clW132bVY8+dz0xbQ5++u02
BqXWSV76SYyXAx58s9jE8/3K5Y4aL6qU6GAGORwBq9Jm5ZDFLg3xNHrP7lUa2YVGxiH2D1Zikksy
nHgI/zmpK7CQZDRknrromdU/qCTbLs/od56Tbm3XGhw9L493WWQ4wsH+zX8wOEwoxwrMmw8Oule6
OhX+GDYrrWpBKIRq3unvzAshRBuSOaGi3NGQuLfWjqNc0a495DJkDJivvZ1kGcddrKbeYQRpP00Q
2cBS0sgQfSDc87uCIUjn/5UVPGkKovTRA7RWJkQZtvvDQYpwMjWgFcNvqgyEu6wcz+g00v67mx/h
d7NYUZeTVKPv5P+338n0uyTZgZD8ljm/xIUQhaHBtHYfwrhuyzqkOftxgWYGATcD6C+xYbvBqQp6
POb3l2pSIZ8GEo46qBw1OKifB5LDauxtVeIV+XMQnYKEVv3LC8mHLXx6q2P2jjVYIl3Hswd0qtQF
LAtZB81HIxdxYWJ6f703jPTMlezx8HHHfBirHUd0Sts+tiRv9iT/il2c7Qm53sUJnUmAsCMfK9Kv
eIdsBg+q0f8tVpF9NBifqHr3pn+vf/h+CH7PwTMtndElm3Mp0YT4lervskbPZwJblM6Q69nUHE7C
6iMc/cpOT0Bc0d9aQBnGVvrmJgJiAuSUaSREx7DchgpW8b2/LqAiE5/xaZVOUFpJ8RjYRuzH9j/t
4OGwlNDlZ+r/VjN1xW8VT+WHRJxUfSRvs9y1AjxbgsUByWlijWhyZqbcZ+BMlS4bmtRZ8eLxq88k
rR5vquyXYGGnWxI33/dPYUscglbFxiN2h+AmIVhH7BcfV1gf1m78Ie1smZ4xDYg4lRbRhVyeOBSN
h9W3Ws6zRZcVYoqAEZ5OThC4Cq6B1M0zluaFsJvSyYgH0cYVUEqdGm0+fZmFuJB39T2LtchBa1L0
ln/4LJDo76gXUdr9Dfyp2W9AeyAHCdwIHoIvpPJ0kE51VowpNLJrwhjQnHEUD1r0L3gR8R0Sm2yj
gVlyvRuM/lGOcwcF6n8oeZlvcv60zouIJx5UsYUVd350DnoriySggvq7BQQXlaGcg9hRnLjzhFsp
eH10PH8EeokRVUl5ZhRharcVltThBBMjcxMvbnhqvEjqSQgaAblwJqpraFm0oyaEaYE063nKBbW7
W3L/s3RrRcIs75fp4anMl7lgtj+gqoeSPMRL3RKsDqq8AK4cHpKnTHp2sM2jS/VFD0N/w53FlTQ+
JBxKGmbElivme59WiBpnjhf8DQrDtbMuOlt0GgkX2tjPBTqfkkacdy4yh++iesTKYP3ZF6bfQx8o
h6pRtUMNQ4gUCC2iD3DiV66bYvaX1IJkYvHeWLrJDLQeoPemuumTSuQymZRQRLUO43u6rU1CxCf/
U7hBj7sn4AwNDshA22DE1VKwF8pPai1K36nvN4Z1APsjtbGfsLk/Mio3xN1zacIrpEWO0V9EmXfR
TJP65D8i58kCJNYilD+Sojavb4MC4e+4cjp82vP9t0/vS02mkO7nw/R6rLbTTAdJIz7W4Z/r3HZc
WTBc93IC/U4rDBB8LUZpwnb5ZtZP0IuucRxje44t/RCMVxqq5X+FedOcpLV5kvHIO25s5zNktVVe
ilMD/yg3b6dwiWMgY3mU+mBJu79nvrjNIcF30OSdlhG8daYdCy9SqjgjGdibPvA5FEl3ljTJ7g0Q
CGCoELsFEjk+cD3kiwNf4pRCrmadNGpNp3qfmTgNpEBDvkBYI0hC97iRqtqY3V8cD4MDKjTEiTlj
/tVqhWbMhXZc+6uwTanb15XxpNxY/QGEtbLedtZTHSMY5/Wo+h6/QAcpDNm2cE5gOfueD0/gelj+
7Q/dCj3RNjjC7guMaHjv4rlmgcgVnV5Deay59MdLAvezacrIsgQshkyneTzg0zkcFCZYyOjCSpmh
mZcSI34Vaak1pdFWDrOQ7suZMtS4XacKsjtTCZMoIReQ7NZHIS969TIjBmm7Kbd5aQaQTEKL/aSN
o2wmnzSbg6C2D6g8vGJizgNp6hz/kdQ6Dpqhg0MeYs21Zm2Oq8f8Yeg91hvyQJInxRtU7Gz/uwRu
ckMkpvGlGIqE1iK857RYZHiGJtGo+ssD2UQPe5UycTKIavPMKQwKk7aKEpCvCj4l2B9FXMxrQ12Q
8XfpomgO5dS5ama5FSgpKB3VOpVfARbrnes+jHkpJqOJgEW7yIr06BHD8wjMWbIbhGWiW46t13Uj
tzEdS4LkqcYN1PkbVbm8k6MjMLz2M4znwa82tCqr2ct42+8ldzWr6LOt0tpJxFs/JYiA5jvVsUX1
u9uBn+XGvI6kX2YJvkPb78lI6HbqkIlfIYdjIjsyPVYbqA5egGN6TEthqKGj+26cK5sG6XK2qFZ5
VjVm0xPOEwf8EI1PjUurabrT0ByHM7PxmH3dF20hVPLZKorj2Tr4baLbVYTEUglSmzHwe6S/j8hE
5s9QuW6GF7MQvnF/fW7BC5lulhbcXuIC8C4QbjEUJ8ddMt26AmaNBbNFzKlEvWtP+mE/s4U1z5dM
cts3EqH9tfSja8j/8gDU1tdLDbn94JSQItjfXR1wZodFfegP7aZjEMFMNw4Jt3tEHgq8f8QsR3Q+
uwZUljVrGhGD2+b3otAUx8Icw+yWQkDKf2BUwo0/F52Lv+RTCxcTvhGoypEAgS5QmkjUHeuup7Wd
K014ojKk4cGQkZimNaywxV3kWBUEJst8HMHhs7zWlRKWo2L5WZeB8CsgYgd9NBY31A4HiraVCL7o
Ua2vwZK/y9tk0FfNo2PbpTSRDn6tiErF/qR5dH5D1Eq5/F+nH4ipTXoMMoTZI2UzUPs5GK4Mvqxt
9T2pGt0C84bLn0a3oN0s2oxiji4JXG5KSwrfH0wJep2pKfCX8amL6tGcnDTOnCl4Y0HJew4q90oV
iTH/l6LwUlCDI/tAcrRL6c3Vi7IryX4rmXTCRBJZcQrVna88xFrm60V8879JKoeDyfnPiVJUtski
A5l8ALeZseV/k+kmroOBCWRkAiHFRf8xV4QXArCfE9IhhQNCNJ+gjw6lX0yiRXYRIiebBTKwHFQ2
PQH/bUHArtu2StZ9gGRmpFlUemBQmCgKnulr3NQtWWc5VHpavIcRCDZviTIfFgUY6Nk+AapT6h9x
jlkdKKlYin9xnTqsQQ/ypH1ohs/sB8t55bAsyBQ/wpaX5HqQ0+sR8QDKcrO/sbsmL7FaBKgbBgR7
G+wNKqnhaZhZtQzqSPZJo2ql3p4AjpzqJ7cw5zYq3fsASYFRsQQGa4iEXDaDdJt88qjKqDa38YF9
z0XSRWkuzh3NLrpImuPBO9JJnU1fW5DORxm7Ovop06zfi4XdiYU8rBFMlpXRKei7BT6MKuaOPZYP
U5LwUgoxjtMDy4OVACdyTACr+eLmC31LZGyJHg4I4tQPwGCwhMBFTyT+B3naLTSSU5vCt8JGG8Fn
KbayROgcmo0kOrOIlMTL/ABPYXc+j1KlBMR+KIftj8nNDPJinfvcSjiRzYPlKpS1tRUq72WrG5Cs
jB9srgRQVeylF8NXjVjouZh5mPkTaEhhOjYjzoxrwKfCRIY3A6lixSXqwRPfnhqcVjd7xaGo66rx
teqptBUQ8nBv9G2uMEkeZNIm0rAvHQrj12mHhNukmiu6lR2/DZBGZst9L8YB35kZkS9mJKU8YfKJ
FX+CcHJY915AXHRSet4bM1IRIeg47Jm8oCMh+X3nwBFGblYNFa1HoAk2h8BNOz28qBLnvt9GZhKk
hpbOnamHk0L3q3fH4/gah0oBPXyL8OfqEcC2s6T+2NouyBzUn6PnQBsGj09kcd5BxVWxHKMQ7Zkc
7LxUnqIu75T3dushNBsLe5AnGBED5kFTQMp/t5hY/tY9YQMURGLbv1/emsYCxj7hunGls4i0khlp
p+K1ImgjILZQPS5S8MvZcdbbHEuq1ZDMs6rPuyPMm4YeSBLbeUV0loF6jI7DpHOyRMkMh9WKA1+N
DYrO4kdBUx4zTjEpU/k1oBn7SvhR8JL9p2Q2MEnr4+EtN4Chq2Jrqq0ztXkEV1bdsSPi6ICKwj2p
WV6ki3ER4SF+J24+mAjXBd83TcfM/Ynmn83FstNA+yHEEv7ECRWemA9ps8NurMFJK470pDmiCiGG
Jds9DFQY2LCxGowFHP5OQE8W7Z4S8cabVuIg9r65SJlMdwkrN4LR4GH8cux9qDQRP8q5JMEwhq2U
zd9CdBwrQodtPqf1eXaSZ0puDAWoD+Bq0CDCMtlpHovC1nwHvREbSeBfCZuDQ3DNr1aZABTLGemG
b5gS2uaGOOHrQjQaQR1Puf3LcSJQxIBntFREuW3HF8LuRajmSGcnSCPSK0YjZ6dXTvOK4SKLfkyj
EdAmx6zQPmkxKTOd4tpuvoXcHquvIAM6umJ2TGtrjy4iDnvOetUIJew0oBRC1fol8s1ishAcKkXV
CtNGFkoGlcAt0/qsdinBg5twMCwKZRvUsZ9Iud/Ln5H1diCbcAaRmqadQstg2Zm275QISyuevpfe
2G8GSjyKjnLj3RKG9YLQ4gi2dBWHokhABpCTnLhD01ma1st+zjOxWi781Fcy8Fe0q64jvxjVQ3Xr
01XWpdr+a+Z9fc0mYsn8G1Qb3BM9KqNOQVtk6CcfFzxAKc3gBYlRfoEmqO6zYfNZgd2iCAzbdqEL
g0uwxdV3uOj4Gvll+Xdg0psmyu7yb3OXEdfm+1zjZIRVCZu3vuQ1xx69GZ/skcDOBaiLGEwlVoWe
gfwaWcyN7e62AfXiDW9/qP68dpz07r0iq6AGewacjYN+Ft3TxDOj61bKQqhSuCDwF5WEuDIpflPz
Q43sV8y5E4a5na54WKWtjlyiB5IWHROZPrbMAJP4Lj0pTwZ2vb10uzjMHT+MuzF6DK3rEWTv2BKx
QXBQByqZyabhdP+blty7EnKeRTidtAFWW7cEy/G2JAAqqsIP7UtbsQNuJyFvb7xLL2qs7lZoYVlF
j7oEtYyNYG93y1BQHc1wloIZssj+gzG1rVyxFL5E8zlryLp6jmQUJZDBnT/o/fUiicNA5VqbK0Nb
9JQOQN0lDk4Nm1kYAWxsb/RwZ6gAcUJQqnGmOqOnSLe3R7RR+QQLmWBaCMA7snSlUjlW7gHzedJw
iWrwsH0ZPM7SjfhvTcNajztDpxK+XJaVNmDCB13D4gTrlxf1glqQLVvGtamBZPweaRWPKrm+JBF6
rOSgG6IdKZgJoDm71cce1+cQAeDzUF/1ec//0WiqXJkSiGGp38pf2u24FzVLckuwve7YiE5YZ5K3
d2CITmWItH+WnskqInwG5I4iH04hT1qiBOVdiko4UyfPCk8VhIwthLH7fXwFG8CnMN9sAaxt2L02
OLj8oQ2EUDivxuDf8DqcKRphEW25SZFWozYDrZ/zQS+N0ooeVMGXh9Q6zpv/7dL4Tagoraozy+gu
/hCeezBPpWMkMf3JNZYPjivRObqXw71HOP9Gjz+WWrOjLTlL3qJ5HhRZ73GVSf81weG3eh8jO8vI
QTlpn5+c0rf0qW3G6pWAzZkafwK95cs31+d+v295rCLXAVYQH1/HTueeh5/7tSK6RHBLFDwT2AU+
fMxJSiDI46NsQFCmJ3xVr2IANOZ64VeBNt3ep/RO4ryjK0lUkpk0APNzChfsPznw+m6Vkm85iINW
fYkEDxzSuUasotQ1fOOOycymgtq1Qj7FYYuZQUaXps7LVDMRCvQlqbwpPhCoa8EXNbdajEUuf9V2
zAilaWIdlqXB6Eiz0xwaj/4pDyNSwac1+jPBXvFeo4K6+Ko8IpeVph0jKYpZEMuuXEpR2XUQgtkW
ezyMQ7VfTQdyw071e2H4g62erTg0WshH59RIMODnk2syfmhYaOEnQalM6loquxOvVjVx5sS0fIWp
fsfR4dBZl8KEaisaD1pHq/QY/prcI9YryuRSh3O98RS/5UdWGKZ7xXUhysbBBkAz8WNHywe+OTDi
9367KQppZnob5Fy7hje1BpiSWtEWSz+3SrydlCoKs8I+vHIMpDb9v+YAsF9N+43UeIJm+rdPEU4d
vB2z1cejk+bOcqRpA4J+yaX2NXhn7N68ELNv+IQ1lY9JC5KtJ+bv/+ZOxPsEkAh3LBfrdHgkolhH
l9YPkLqsfLC3l7o/lPNRBLod+jlEh33k04vG1dp9htxq65gvAC3no+pZvq1/j2Jsl7WgesESlUtX
raAI+Uw6VNReNs6iAHYB3vLcShecmvRgxO8UAx5djCJui/soSNors7W6Coy1UUuGQ069e+8KUSpr
tXCUQWjlL8GPyITZ2yBEEFxxTKYQ7CcmuC7DYfp5Ev2qjQYU/kLxH2aPN/PDrKsVanXDMao9L16h
fC1EoAyDrCAXeMa5J87DU8JSnnPT9kW1g+oBg9IxtPrp0DaFB1mMXdeZZcB8kahmiEDENJSZ7Bel
JgSYOCdPrXy4cqd12BFP9hjJVMSJU0YqU0gR9DkCeq9xCc257gL9Q0E2bo4dPh372cNNT2BVfebY
9STa4PjcM2hVY8PpCCfGwU+P0B953bl9TqnFJqgaM2bmgwWPikkdNNkW2CAv8p88TzzcItyex8Ad
EbZcrnLOTqH32/nyIp8JzQRGCG3xM71tLmNkmXsNObF0ig8OU1FmBgV8/XalR0lSbsZBVvOs6oQ1
EEzxWxUlFBZs9cBp6266URtk5F7KsoqLFkhk/x2ssrVbgAO1xVaXWwh5tnaNNYh9T2dZRenJBD3S
8iox3SO+CK/umVgoetYnedGChQsrfMWqx2VQ33gL9a+E+39GQfBcUF+zA5nhPiy84i8qhLkXBaxf
25MrSyV2XVQ2Y3xWIatSHMsLCsoNr2/DPDlsDMYHlZAgBH44Q6c+6fahp8VykM1qBXyJM1lRBsNp
4USmuVCzBSU9rcfdrFCV4kj7RMqU1puh+4VUP6ps1IVf337FJaQ0/UbDgdpku6rbhllquJRSuJPW
OaaVDfAdvmyMjk5y7MCKaMob+wh/DplGJf9O5XtWDPBgMhpqdncduj0Vgp7AFPqVRsv+GNqHO7sU
E4ymQHCOb75ZON6TKWUne109JUfbVOBwrQ4O3b3lw/uAb1w/h7mccBOkHq27RFj0XwwR41iRtyzO
wWTq2REGcbYjgHSqfAvgLURoELnfnS7P2KBMNjQNtMsXtMMcvEwbSjBRvkdn7eO8EyrrTX3sHd8M
vtlQOAfhwmJSflVO5qNRklrh5NVrBv/84pOjYRLQdDOXDM1pYF9I73Ar013nxpDA4q3gKK9L5nDH
TZLZUjN5VJBilBJjZ+SIS04ZgH82u0g7Pk0wkLMlyZlDWJDHVxGH0HiT5fpgFwujQ3juGJ6jqom3
OioAtR18F6DvR5KFux5mmbrmdHGccBUPjjPpZVjZnKvee7e0QxIam1002jqXEZ0Rcp1h1wRTmYgp
vTuplBmnSWxiVFBrcNNTMgWNr/A2nEe8JNT4dkAVe0x7SfVbFmkv/qH1rzvkJEFX7BpbUaxLAj46
l0DEzgtfT8EtvSiTHQooEDFgEzRyFc4iDWLRvIq6q8r8ESFkoc1zWvAC2+Wm9lM+06K4yu0LSh3I
WDkXTLGey2yWuWNkldIHEomkC1S0cUfe+I95VYS8pYAmROHELVmBe/yneNhIVlc0qihGjfv4omfS
Fd30GKXXwxKhUjn6Yq3P9AC+NCdE4/fhQgcSN7UCuwiGo9k1ijX9eOpSlk8lV47Ug1F1GliEBCFd
NqABek7jARx5Dp7BC62bCLAYpGMC1mH753XY8Mz/TWVg1a2NsX7Z5lsqKccTFmtY74raHHMVelVf
b1bvZgiQ3v0Bitm/VGuUdGZQPtlZ4eIm1nxlkNFwxc80CzgO122bmogymzP9Lfmoi7Z9p8qE10wj
auVwPyNQTgCWaYAukm4BM01Dz7POXuONnrjYf5d36O6t8AhvMTj5Q4MzACgVbjx3oCgkuc3QfBWY
xk5U3y+GFsu7r8T8g7cfAqHWSK668CwMS9UwMuag/wvdlsNu/73I0ilxTeEGVDln3YXWUcU+QZTG
LSnOr2Q+0h+tA2ta+9kFweAbUcfnR869CHdsSDCfL0j4ivNiAiy/6Hy4VRznoKjI7xUtub7CvwkX
5s/IHVB8MIDLR+TtuNBe/Ti24qb0872jpZ23wTVX68mqRT4nczTNM1NIDPU4V3LeIuQ/ngP8pvn+
3uYf1Kii2q3kbWWWprreHsn/OpSZ0PUMwgsOmOl65NueekkitcqO5Ax5qsoDJyroQfO9Q6aOktvy
HMimpVgtBtNYu0nbmOdJ6LnbMBMQ1WmvohkesRSiOyFGW2BhEyxWop94qh3O5q9PYyE2i0zP+R9y
/f2dV8rAFzkllR8dzrBzSbEONc/1/noeySBag/XCbtbeSI2TNHDjWB/0sO4mC9jkt6Z5Liuzyvv7
36twomUNacSbOY+yunU76LGIuSdC/hC27BardYvk0Rz1hgnsaBTjv+DI6eKIkkVvFGJ7kiETigEq
pOqn4c4g494FYaEBM3yKqHDxdmOcjW/9+7RPlmNGoDkf8gfxi51tK+i3T7cqcbHdkyS7RUOGRzKf
6kjOJsj1xbogsLPaGWQwPl2R0op8BhwaNqAGCmf8nFbozSkipjpaVyiDvoXtFQWs3iHixZFUfpD/
hOafqFuWzfPwhgy/y8R7X6DMJr/cugpxFaKHzQyeB9yVFCxZ16dHBq0zYEdrhduXlAkKQcttTzbJ
zhTyMkzt2qxiAfUpBF0QbJ7/2vd2muA/vjKPSSAel376+FlEtw9w8rC1J5Hecmk9ClQZ1JDQfaB8
knunnkXHEMJuEGfkjXSdApFNAEaeDVxPhGWX40TsKfISac3gTP7lkYjMMCa1KFN9n4BeeeCgMNl9
W9SaZms0xHrK6tRCpu7FNm90wlt/x3/kvUih9QCcRJB/tIb8jX8jdaOQm05srRklYTTxoBA+E6lF
8fWIvlFNyl1CNWtliJKNw4FiQibKzfht9Hsa2uNwo+Yv/Bs6NCmNqvMGOsh1Fdkro4isIztcKuOG
+K0oM5FiK1H3VXgmylElO3mYKcAyipdL7htC8rSjRvmftdU8smARbZs8m2q3PoB3K50TNgRKC7Y9
kyXj88G3j2cOgGWfPQSJuBSvZfkR4AqFaUgUG7qZjp2QqF56zEjlW7/uqoNCooB23G7qbP32OhJM
Oq7K3ZthVs27V5inZXgkIYlY+5Yzx7n48nTdUgOIk3EX6Dq5EbR/MsXiUdoBBCOA/skBQ44EAusw
IjHEY6VxYjM+B1Zf2imYs+vISm/J6aLXPMEBL6XueUJNWa8/LMilCBXTN7Ml4xr85yua3ix7X3Fl
P5JOvXX+uc9k4n43iUC9yh0DUF8kuWevxecZfRoB7l1NptmtpK6XrNMN6ocX/mN34cx/2RlC5/nv
fWno3FnVW4/tB9JygLCG+8xDRMc5vXiNcXb3LoOdUWYFlimlvFTzwKYF5i8dlKsWrZJfSwgFJw8f
h/Iy5yU7IZdQyqQl4/dFVqkflj9TpjbRrf736LA0a/i9YPHtv+Svz4k3+Og1Pnype+/nZI0AN+p7
sTrpowlGUR7+hi2N5bqi2IvvFDnb7O+J7sMW359hTd9aH6Yxop4dPpK9J2+2IH+KUE2h9W1b+e62
Pr9nfhblqQTviQ6uT6ea2JrD+AKvHzdZ6xH+FX9SBXMS2mJ9Ri0G6UgcC8V7pDuhstWBzmRh2Hwj
wUUG5kn2nUrjoncmG3bfEHbP5hwHk72Glp8qX7MihSpzO766XuTp/pZfJ09BP0E2GpVm/eM1MNlB
hwEFzJZMWARsBPV6bevqBDDRxlKZtKJuLTNr3todD23VHYADZUCt/bR9RbEyJN3NSAU8ijhPMTc+
cM8Gz3who1hOhbIQxm0aM+fUtj+vQRgrG0v7IezmQXygjENqBFjOcSKUcagrGZVIR3GLokrXy0sG
wisrVSnwTkFXq4+HZPBGBypH0ZuCurQKnRVwjWLkaTVUzQcwNmL8QjnstwUP1mB9LVz8VyQ66PWk
v226nPS+Fx/7No/PUK24X/ksF3lgOTuyjXDgX9eaarlFkHPh0dSMYk6HaZaWZJ82SHtzccxhGD71
auPS4vgF+Vm4vyO59nkXcursLOtjiVj9kto2iDT02c0nsGl5HI2tteAYP3f9Sk5+5vAfeuE8ahwM
NMXMEh7TvFi9z19/yBabQT7fYKbfezUJ1IbGTi3H/RnYkE46Jnk1McWfBjS/0j96fA6g7zy2yFdG
iEhmSrkxEvCBx8uSsDGhPs+GcjF9G9yZ0ZSfL6lZKh1HE6KyiU3gFqI9d6vYgc0TzKy0JLNEfhm4
4EQ7enyQPG8GwZ25YEyWB6vnvmScygXzqLZt3rQAbeW3ApAp8i79tvB9vK4wD8TP7Ii+qmfaahT0
fPJxkHj02ISheZ+wFZE23kq40UVZ8j+B4nlqAqvELtNmeN+DtYnqboeG4DLtA7jqr/HbV8sVRa9u
H2ZEhv/y6EHHKNzAYfMy1iFiW/7Ng4a6l7Z+vjbbhb6tSZ2+RmxQoD0SkmwNyGdfr8shxgLpxdRR
eaw0SQ7Se7pcf+nDNwb9etLtG77Ecg1GQ0EI6gfjvCTya/muXM7eoZ2GWsd5jna2nnTGeMXk6Y+T
7rb+u8SUVX5gIqzxYit0bIrdfNZ12kLE4yEK5doUfsn8Pyg62YxpOvgE7lWjFLocU1NcNcj6kp5K
8PRVimMgBYUUzm6+Cpj8evQXCtQZClNWZqdCCelNeWO57CSKgXghJ6r6BCUWr4X5VUlosQs0WLXW
v2D5b7dWqbluRnEHaXs+Kr0O6au1hvsutRmp+BDHi0M/BarHu0thz4783nYNWH7ikxGWWxKhQeWk
ErV/Ormzbbp7oMe8Yxfh5hZf3x+g1P0EcjMWHGm+z87CKiHGJWRdPz72gd9AaX3EjNr6fdXLDzcx
epZmofhvDS9Ayp85YV02eJsA077WeppC3FHyTsUmVFlwLWVEedDxa67QRr4rlzMFDsdpk5dmfU1n
amvQwXKYsimEgt39GpTx50EKVmS0HUDT1CFVfqQyIU1g04fWbMg88bADf8FBq5cSkvmOszJl3l6g
X8wFgSUjY306/QZEhM2ST49D5/7hZPbwU4MYXAuavHrFQqYk3sGH1GMFC1zM9HbndvDlbhG5tKrV
2PmdOwSHbZAsooqW/XsNwdEhlsKm6VwP3Xa6JfcLcF3eE4PXBqFM608/bWSxH0AYv5VgiZzw1+Qy
a605TNJr/c6GJjckerjYsZgQBJ/jqdPi5/kswjKtiGQDMY/sdDowF2Lgm3TXsKKAqHje6dDFOaD4
a+5Th7nL211iTkZTLY68w9x2wzOH0MT/a1ex2Bq9XiSSXal4ZNf3wuEy3HxOO2CEV+yUpb170hhE
yZQT0L8L9umGCqEaf5ZBnb/6Mu1QDWzP0M+R8Lt7WcmwEYfZNC/YphTcFLNjmp8wognoV+6ODGV/
gzj9rRhwimQDiQYmEZ4OY1zwbP3FR+8MzpLozsu/g5VWwWRzad/7zvVzjFTaomE0tX6i/qT+J3WB
SUnJtn1uBWvtrwwessj9vEfDawTaJOoIEZGecQ1s15k7AzWtheOE9IYbSiLfMeVCSRhBhQa9ncFh
Mj/MSBVVZfQh4hYjRpgVLGNm1wC97TGhPjKX5FfALLYAq41Jh1LirfealYj2v9XwteE6XKGrpCTL
UTzwoAiMgDMXjlPbDtbfjG45EBlscBPN8AdpYwF2Cy2R+nqvj1juKAfHF+cfZQ6q8EovNgyEXE1W
fimdD3zniarnHcriFYj7yFcQnkG77DtqIFRYstuAOCGwqLb+prhuWakQDQxaKlP58RugNQEKOBPp
fyU6vcpuh3TmoJAK3bCGoi3DWYOnjVU+UBhPMXIAhVNlUxxzAYnNKq6cWGh4HEHKSOUr9Etm7ll2
p7UnkTZvuU8+V+hQg44orpdv/1pyNdTuaZySYCU2TpqT9Y0ByqZCo6H919nQVgJHUt5SfgyQT7lG
S9RnJ5ERGQSi1FTXnxWh15Um6KaaYmC5wGokjdDnOEpxaV2la8UD9dUba7+aKptWm7bH4BcvdafU
VzgIRXYIRnDdF5EpOw3BkSdk8juWXaB7OqTNBABpiPpLhr4jg/csqV+nEllLp81vFH576dYPHBW3
RdbQIWIAJsFTscrOIIeMeqvPEKOqLjpmzhKjBC89e3C6j+I6qplNVIdIzitS9jGyZ7fkd8lhZUSO
1COpLw8JZK/e3PvaBk6IOpsgoRvEWEi0GkONUDN/48RQdECUkapdUCVwXtMcbwyd7mnoO6/1Sp7D
VI8d1apKZgsN6zV3rX3NR2xmqLQ+xyqpStZZt1PhlHRrItirS7AzyEFfsh7rQJV2KB5aOB4le7gL
Ed8vKr0ec78E8ky/TJ1tMT3kon1znjH1qlRADdL371ssQjl4pO6ld8WHxrooRmH1VohsoGyOFg/T
IZe+9tF6SGANKK1sHRF1PmeAzXFj23w2Amjw8dG2rsZ/iIKTKBYuyeHbK0tVhEoNpSZH310f3N+R
+jBJUq15ntfanumGcHZy+tDKkLPbW3eZqaCEbmSxkxIb5IBCHxp4BKgkYY1EDoBTA6+pEkjXdnwy
reubv/WNtOVZZ+TTQ0KEtNlfhpOqXSxMrjBuvr30TS5HWgnnomta2BeGKA+c3EnYGp2mLN5QVx2y
CvMCN+cONFF39LGyXADSXxpATPIR7S4H2psH/0wojZ58gch3rUwQD05HgeDnVoHjTS/zNX/4446u
GZBVjux4MmDCPV6Sdj9v1GHQr8gCk+v3ZkGvA4VLHOShq0Qv9AsVH5eNRi3eekJt14yhLN948EJO
d8WDduCfcoaSyjASFWHsvnyKTIek1HkcHMVLuNS3o5CXR7SQzGse+h65kVL3ZQJfcuMj9E/TDZe1
Vwc53xexEsKlsvDyQv9tgSYMEATS6RVX2cdSjn9BzFzbGncGYG4VW9jNJ/0f9Fpd2vCYpj++hrD5
jrwIHIkhEiZkeNyABs4CwOZIXlrLKfeeXN0luRd6/EDkwqg7s7QbZxpElMgsoYKwSJxSf77xUJZA
SNy8CPulRSOFon416pKQY40oiFCaYIBIi8yB6apK17KfCLHI5hkj+VpmlAQ7wcHOOmqOSy2iStPb
VbnuidGK8jSu757hUPF920PVN3l9W9wajHBcoARFM2PA33fd/IhgwNwuGjfWTWLYWBM6iK+W7J+Q
mVEag6h+5uFmGeI/7pylZqMbejIopYCEfRSUhvKbklLdmqkGQwQNcDfjpt7vlNj+RcVsYaj3dPpD
/ce/dLUbVaZla/djrTelA7ZnRuX/ae0jOvz1JuQ0hYi5HjJGMwTdB6pJMqW5hMpT8/jXax+QZhrF
MFEtR7KaQFHv04LmGW+/yZDFqsOnJDRu91kQj9JYx1gRb2ps/crbBdF0lcq21p5fjQI6JLyqotSo
Z9xGDUp2Mp19QmgFIPz5eVxvJ9RsklUgvXSG/vhth4eogHlay51hZ+d+SwRgM8H65EP/4IUg4M3G
VaJ8ItJ//ARQu7B0de/2yIplWvqCF88Po83KKHwgTstyXNyguccXCpDtkU3uEkDJr0BimVhEHPDa
TeFOLepwdcfGD6Rwen11kyO6RzZ+AUpGBIy/1N82DoeLqTciGb6CCKdb+6W5mhYzBM1KoAdHbvUY
BrvtEaGjUnYoEsbKrmAHIIVMHZDYlcwdQgxoiWwwn7D5Z9PaW6pGpkqaB2YJrxP9GHE7QgtxPVhl
77Vkr7uW3l6+B/d+OaDpBT1Ugdx64OZR78AgHQvTIOAxehULrVZb7uPliQfR5mmaNCVfBmMu4rhs
yudaTO4py/FwlwAJbCnBpwMlBgfICMxAO8gLP2cxn6dR0mzP6vsI2H+cD3S99ITOIhbHOFT8wTMm
/fS3tsseeyVckfEkGFRHaFxcNAFH6JrJ1j7Qw7SlMoBx5SrZYKCm9/qZNq7JcvTRV0W7TSU+vOwh
NcJPPu6tCg78YLJAvWSfaprVQJWIHVHYge84PlTntOoDAwlgLvZQPAreUfxVijrjulJorxMRFaY+
qMNXMmuzF7Uc9wboPgHSw8AgCaymWD2hNCplnwbzvEIG3ZWI+P+JJQ6MlLISG7uTJIKwsneANMJM
BA/SQWR7XV6cn1wphxuDLDO9aPzzU8kQkxad7fNsOcO/Mw9h859NURd9BURF6aP/Fh6Fz7Fuqp5A
3Oqwnew2iZNzvdtu28npyVTzZkdU1zkPaYP5AGx9TZwYWWqInw+tYnsGfbmGwLWI1hc2pPuRB1bN
p7UH1rVZmYjcCZM8LLZoMTqgr5N36pe5E5W9TrVJyW1fvpyWkAvJES7oKxRbB4q00ZRZ2ephQalM
gXZGnmJc03KXC7bUdMXoLDOcWEpqIz9Ab5u0HrfdSTARvZfjO3B/BJFJ/vzC6cifcEuJ9kskpz7g
IZvXn+YYmHIz+WxQT0Ahqr/oE/FrAh+VFdxFVYFE75Plul44P7REugzCzStWrZR6+cHctSCnRssW
aJX1AhlguOfvPl2g62vpTbUEZQyTqZ9cxpQvw47VKtuZBs82kt375yERK0eK4IquQyEyBCfgjSYk
FV8wJTpYjp/LfxhueFWJASHZlXetnoN/M+a4bPRCyTnEeG0gB5fqxegGgIIL/29QjKWnAQ2kUVvC
Gb/TUm1EOhOxPvQXDXacZysz5bHaS4funV0xEFE7pnZBC39gxE+0W8tkBmW6Xmxq1xyXSdI51qKH
cQjPIn831FpNJBxhEUBefzQ6oLESPbp5ekjkVEsHoPPXJLaqGLIuASwTNZlkPriRLvfaWwqxgIMp
p0NW5hSMNpozgI/hCWugzRQR8bfstCFVmSmUHWCOxn8HXeOFwNGeGPfYVbp0RjESyW12ZqmI7LlK
alHNUZRf5fOhDB9xPgJDTJwSQxkg/gW1YgSEH8oD9LA6V7qo7xnDH+S859FlaoGoHq4ApGZm+Ls7
XqLm9INRhZ1jD3JjmEplUiQpG4RDsHTmzRtdmJXoNlInJmxLIXLgVUwnhLQqV9k8KIhGzI/QeRkp
YXaTb2vJ7tS5bEuHIxyvwOdymajOCKqMuYRywwyyx3K0BoifJrBaoucG/Tdbk5j0B0S33IVQE/0j
eVGC0ycXKJveOZ5j0MzWCZPh2+kAKP6HONH98TWduKaxZFYtdbLCNuriZaYftJsefoo7ihxcUsrU
x7UtBxIEr51XrA52/2aIAVv6VD2+pjttq8c6BjLld/5rxOFQiWXM/RsBww5FSRFw8Le/4Z8zIQIu
wYIbKKWv9UlbISCAfTLc8vLRhxwAk0khtvOQo5eQSrE7eoLENmacuxGDa9wrkwsQYnyJd+WJ59Ii
xmmOtUiTZvbmDXuumuhU751Xf9fLXOZy3blnfGTWpFmeZSfuu2BK4A3cponw4vPpey2+tEQPjLZN
Jl7SZ4yiw1qTfFid6iCZOpmJvGJKjyWe3KGgPrStBYt6yzQU8XcS+a6zlsgcRJCCEBO7Wut0qIWP
aG489QxHqXJKodZ+ur+K7ZqQlsBE5/8RUitajksQpveMC7zZXqvWfE6rviCnUOMDvVDKdNdgD6Wt
ljwhXYsSoD/zSCwuwv6DovXgnpZ6nusF3KQtdAM+4KEEZ8XOatuBH3qaJDgAzvahcbBJhg0fazK7
nzmHie+tSDnJV18gji8JGAtWt7Q3fd43p5BytYoajbwkFjxra4D0dRABZ23V27PHNuVHq0WaNdxm
6Z5OHPnd/BXfAHgnqYeroxc31weAN3rglu9MmNL0FZzeNNidxN9UWOtbn/XP/+azPJQTILlIlEu1
okiTZVas5a9YxTzqH8wTfz49LG+wR9X+V6CuCH/Br5MOfW5QSSUqIH5D2YSo1iSxWoxZPkv3kCsQ
6cClF5WPue0v7G7UrMAC2OKgeKzLwEfdpfmfr1vdwyU7VYqKtPYkNLelvBf42LFjnDF8nfI0VsDm
W04MpZ9Kzt3vfMdr6BVM1n3q8vopjQWeD6cl4bAu6pvuwziLEJIdxOKZqNIDuf0ci70KM39e6DB9
l8ObHRvQll2oAsMMU9pzftifQWV08syovGI14hUE+CEv9qU+WfVQUHaYJsHRJW9ftG47bkUJOvFp
QCtVaoDsZqn2YsZSVnEMiJDh9p2RNHrfXiWaMskNVMzwr2j7y8oQO59nRIMLkR+LaYGRXbK9bIrR
+pPtjqrkIav4AWLUH9R5Xd1PHfX3rjXaydSzeykUzVUB4boDKfVZXwr5epdxbSyZ/pnhZdEw1mM4
KdwANFZEOlAJr1MsM1HVpZT0Jw2XJDMbHDGxbOw6U4/7w7zKa/CZ5gPz2yc+AfoLr1TZjiPl3SrO
wTuVkvoeIHQQdzQQAFFtDOnG7huF4T6CgTsNtBA6OcphpCx0X+gpTVqGDHD5ghpMuB5laOhGK0Nc
FHfhrQvEvXi/UFj5/56eIUZd/4loeLH8gkcxdDEHA5bFHRDW2MWWTg8K9SzM1WNtaiz36uaiYEgb
jxMJXRrPnj2pvF1ESgeqKkaFVWJu+AGvtXa7AtVgCE5SF8wc9e1N8okX9yiBkL/Ozt7OZ5YOT5Sm
Ctna441dlo+CJZfJI84SnWNIPSihNW3Ka5ZkM6I7FGFaxEXjyXegeRPsWHtl7RGOfroGUCpG5ciS
ix/mTvSLxYGZYHMl/6g3F0SFpYUFeT7hP7M0radzbHRKRsbkZs+w1DqFc1z/q1nyxlMX+GQ9ihII
Oz214lMaevvLSFXo5siELFSPdNz91Wo6BptfSIafxeq+d8RuZ9h4xEfCF/h5a6eDC9uILlKVnbXP
tsnMhjBiU32V+UB4buuzxSwmb+ZZtdnN/zVww6tLf5h2CNKTHx3/GlHv1E2RWkLbGoDSkPHjlfoI
+F6nx9EmWdMpZ5xP/w8OZs0d1E9MPZ39ruVH33SXp/62ZoCgQwq8BwzSCd074fDziHugk4cfSoZn
/OYJJvy7JMAkeGyIAt/oAFVLevwLnjkdA8+Zlv5lzA2iBxxaAbkb8utDedihuLVEeElK1npMXgwB
4XjiYdrqVdhIM/7KxMB4dqVuXqyLi/TPWuanutRP3gwEwOqJCfdpit4l8mrqVl7F8G7zzzu+FTfk
U3AWUcIUwdYsIOxvaaxt82RI2c95Fk1kfJhUat4uihrbslF/57Vodv0GSWh0HHXXG2QtnuovsshV
mPBF7I6vrfui79JK0gbTOURhpVut/Zj3jUxJ9TSR5QN/rScpDek4IadBNwlfrZv0iOMxREMOkqLc
WAqrx/EoY8lBzYIFKCDC7VAXTIEWkCyp7BhGCbNhsQBdWO098pIc/CcWTD7n8IOm1aUTQtywM6FZ
gropVB7qR1Qg8uZAd5oxN0Xcagq17slKhOWbUFDo2pJTz0l6dhZ9dzoqsG7EctjsrVIkY84RADPc
tmAtdMef4vkZTP2EMf+R6QYkSVZU1lL6BK0yCrMPD2GFDOH0MuXunYYOxfo/9C9773XweT49Ftz4
2soVSrZxDgGV5TcJLyyXZFC+2iTckym4EfIx89J71BFAPCS0ZqxL9kgtqFcOgFwoMWoG01KwKbG/
vpFTOQPjzPQClOgGSCCk4pCbj5JFjA4NQnXL0GZ87MnAZMmkv0ZODXzgNpLTXhse/FH2CHMPQHjj
XsZBDQFGwF+kagj97jyD5/WL8d/7Z17Z5Q6gKzDEmRHY7KB8K+25MKBHqcDmY8DaLe/WyUhcYFtH
crLlj+6PuYElf+J3uviFb5e6qI41bkvmVwtg0XRlDMlCsKuy5MrdI4auhvCajKz9PLM5nIzx2sB+
LGN4ujihRlkqaSR23SZ1Abx2Up1J6FSR8etp/r4nm/CjjTkd7gpObnQgFg4krsNWgp6Ll7VIghIO
cwE+KMdloFQEsyHcw7OIVibVmwvvlWsT7vlootePrwCZ2flTDCaFes1e1HVxpR2s36Fp8MGQKNWI
wMYdz3yeRqdcSy48+SnVPUoOsSkbemOpOqBNlWObm2F/Dxj2N/TZrYlyhM4sRoyMbtEsBXg0k/B2
yqZL4wYkzGDp6KSaL6x9B38qJMCRqT/R+hcgQbmJHlKWQewrs6K/ITSnbMaCdZrGjTdGMdCbqQiI
d9bNqCBKEgl3LcU+E6gNa41WsDxqpWpmMiQ1kUsTOE9n//MWJCbOqr2lkEPLyyV2Zle2TOpavMg6
tpdufRwnfYax9/66+poyEYXgUhqqeH0H2e0SLZFZ7UTDQgau6OFNVbXY+9/UgQkECSB/Gvb/ODRa
PZ7K8RWFuSPACwHsohTmx4qnLcjOlxnY8afI+ewfqV/eO5Vieuu1wX2B+l0gO09SmOYKvSZw7/X6
dwPGDUNIsehIryFd4xEhu4M3zqzh0TyVJqfOphZbUnZSOnRwKsCblXP6i4rg7o5pEtI6tOSvn6C9
ta0M9D/QPMWA7sfjlRGVxIahlB+AMm3/EHy4stfPcLnXzwxnLpitT8nrkPslpwx97Vn21RSgdN2y
K0klCAI3RSlEY9UNZP7NEWW9/NvJpsq7PZ1iyrAGASR0qd161Poruv32+OkU3aNaHEP3Mz/aOtC3
t4S8IHS8eMyfF2fYnKSSISLgInlMbHYhuiny7VLFByOehd5HJ/Z/GcVK+34Yyu1CKQ5soNJvyL9e
D4nidk5HHf7GGyBnfUq/keCt3Z3YN+7ww6x6QFCUQwd4K4JHzk9B2Z7a9+wCMWJju13rr4llfuKC
LHxqxHXLHQgRUKwyWzfJ01+WSZiAn9r+TcuJTsaMdClaGl49tG8cMsKz8PNeN1VJiB/4DTwZzEj+
ypSW5KRKxvAGQJ54HfYWzN13EL0bRZI7sAXwY2uD/fADfc8IvLgfvuuj9tTSpwTm/SfsK9APMvWy
YtncQ7MlIWGTYMGdD/p2k4VjmqTTy5NblTu2Q09oJ6r62hq9+OiX4+n3tDRHygeyproAma6eiFg1
gPFNvQBuVUlHbipmDyEbZSPTH8D4g1iEah7+zqqFcfcTTwzqszDBqQY4QoW1hlAYLXC0GYlLBYrx
MTBpg1ERbTgP2rGYxiNS+9i3ptoQS6OTXymyUSNx3NTv46VVT5qb1sYf05BecHme1OJHYZdrGmJg
l2Jd4z9zFgrbRYMlbWkBIbKkI/juIbopoy8ka4VJG2VAKDHgHkmArW+5pKqF4nn+mAOW9E6IkT9c
CY1hCvs4eMtE5EYIt8r+Pbi/yAcaFGIal0mlSdQ8ioV548EBTk3ngHn+aAdBXCL9rxZpm+F8RPfB
k2V7/owm/vp+9YdHPsQNXOTnaTR71woMBMD31hRchr0WN7IhGczJcr9aZRXsCleHlNz2y93CKYzc
3ZZXfJRr90b3g4QfZHl+ONUGJD9lpHA5E7kj+pqPL9fp0w9i+7ZulcTs919jJTjtQPcJc7DDanU5
b0hld0m2fArxGrosTC8gK7N7wS1sSu2+irLQWFaNjHtddT4l5cHa6x5WOjc5SPZ6ZPCROF9RJ1x1
kdKG+wr/sgr0yi4kFyCEPTf3z+itfNd5uwD9Lvxvk7gkWYgojKzcc2WagbtSCFnziceUZFNWAS86
4Hlw6WEV0xOWI4DX65NGjTnYxUFZ+KgrsEEspZFOuOQ5ecwqEzyfzNv7hnCn+CKInjpc/MrcFsj8
7kuZDHk+6RpgDTqNsjrhUB9qvFRLYZSKp85YZOYF2ggIpfKAUHWn6NupDVuTY2vGwU3NlUA2uu8p
Nlw33Udj0VuenfiKsztIPqTnE8nfNvCLbQBVHRBpmzCfxunm8+vvr3CSFjngxPDNK2eWFviRZWf3
H8X6+1cxvnUp8CldZ6eBhGveDAba9a5tvMjfKn2uLtPfiFqhy648+Lhqehx5WDsbyuupp3oDj+tl
A1wvS98LfCRejh3jEQz1NDCn5iSzX7WYW7MqUgEAZVGIHC0M7Ahz9WQv374xSBctd0AEwjATMSEs
X+QwV4pjhWijSLTKxXXDM86jn+ExCD8Mn2z7JaSZHCl9YB/UReG7T7iNp3RpyyM5r7o3Vqj5wGkQ
yqg8l78U8BhekUmCpVouIr4Gucu5VLQpKRstnI/wsXclVQ0bHBmjOcmx/1QGo2DinEtNtzzPVxYE
KB99r1623YCOyQ6N8f8JkqYLZTCNh3Utj5UXpSPNIXiXaVIwRxaOEZ8DETg4DEtJgS6DFf6Oyi95
wySH/g0K78LECzI0T5dRBoTr9i7H8l1qQQr3BcRILmiqgPGA8+ZltTGcQVl2e15W1EFB4BzEwZ2z
OOAbbVsMuOkaxdwlWWi/IirLnzc1G5GBAQrHDLezpmMEAsDmM7vcNV7QuBXOcuHpiayK3tETjqnG
8t7FEGg08QK0Ka1i/sa+KEkqvcT20fvMAwg62pYoYd6hk98SMBc5g/Kj2NbSiOhaOIprhrrGrHic
7ARY4avk/zwl1YoR0MxYbviLNQcMl84pxpbWyNnN/LxfqCl3ym+IMsBs8PdYAkrc1WUCAM2RNjlP
MVr8qzyLE3zauOHzhHJQHPff1dWobpTV1+0W3SLzfzNtUDZCUrrp4dAxVlgk9OdJxOOpWcDKQkhM
wDQe6ylzLuZOco5LFxdo6jQAEM5HAPPskzeVg5G3GULi4iP03ZUr44Al78Pk7SdOS1cRAkVaRCs1
NJ8XmWXm4fZtsnZc258ChAmjaY6faxYDkA2E8AYpyYUTrNd3DE2lrT6qJ8vsM5HHPHBLqyqm5OoQ
Wczlb4awziPFh+i+caPSBTB/H0mXVOlokAxSq2el07GRRn+w1SbCqlwURqe+ILMrHGwvW2NgHxvs
gyIISO4bIwM8LNO1d1nVri1lLDDpb8hGb6X3spSc2nMrAKjHtuUPSuLRuNAobfQMtvnGWUNOU9eY
+5uzOKihtoZnMrKmkLsVlAx07iHJ3TAdDMWjpn/x3iXLBdmn7TUJd9nAzPvDw2Kd40qLMGr/9ZLO
oFI9KyeWA38flnfujURC01BS0ZB1ellfU2x9KDLsyn5McCNj4+7nGQRoqprATDHT3kb10GiGLrxG
umcYT9B7o3cJdcWQ3FDPwWpSrqT9F+CF0J1FgmCNsut+fFL98sz1bHhLNn3TuObGHjL43NWDHa7y
q87R5pW9ZWW62Cwi9/F3Iz19fIMjGCO89vq2UjYottsqeCWvFEXSW3OEmKnRrrliiSxU/yqYgZNu
sHEBzdq6vmH8egSAmc1wX7axXmY+Ff4mtCa9t4n0AFNIVSTd3NvkgkpoLDn/xOjJwf7yeHTP0Uvc
5kzCcQu5+Hf0R/xrXBrHSbPUkBXpygRijpctCABpAnsxoJSzMM4MlzQdA2C/oXQRxE4N7Nq0V+kJ
NocWD6iHauvgEZCvOPwON2KfHDUFDaTN3TskuIBZdSqM3RIHFnFnW7d8M/2uoReWw4t/7W/sLnro
rtZ2OZm1V4nvcCtxWGNrGz4G+H+4rETbb63v7ZeoIuAliH9jdKIirYC80kZWKUPN46lz/6AF9QYI
QXekUhMXRYasJt9s353Vc3Rfo0XXesXEHEYc01cM/B/tNySAxsyZtffIMuTFJK/0yR2SoB26+27p
2cdriMkjyX/w3JVMNdTo5qpek5Ig0Y1xSPqFQgjyqqkL0XpYdilhLDSsNIReuSxNPEjqKstKVo/u
pxZddagu4s5bvtpfw7NH4qQNx8CLh7vEoXhw2km2VYgMbyzXP09+gYZkIIT6vmtqYYMWZg7pzawR
A0ti+2D6wUR/CZzset0sV5LLcptmag6eZePjCfni1PEbW0urwGojOctxNBTTWLy+tn7EYf0qUuiI
HWhDeVD5DsCuWXniAI0GV/JIqoXIhf0zrOFBkRLj4r4BDfZxJ92hAGjY/TRen7PRwJT6TYx1rwDW
t7lOYf8ETMHgIDwPQKNDPY55LBKpAEYNK3WSRGaWqn7P3ba69B6E5Oy1lOvlKRFs3lQKwY7d1E6E
ALd03eq0hyV/DGl78DT+i5SEhofbg/svszMtWnSwPHyoXNqwyQgnYabaoI+BFH6H7UbD1gNMmxkS
rZ4JGubtQIfiqybZKrTkxidGo+Yy0qU6mYahkcNMZe67186M/Nk8ZCKeAl7nscuMOOhCGP12zYPO
43F2NcwnJz97HDuUjphCWhJ4MmwFiRPQ5RQKq8RfHvrJfU/INFsDo8EZ10GEa/97k8uBNTR90B1o
UVy8Ir+ahj5qj1pGNIv03lI9ZGAdlbNxYyZSlRqBkgfLlBmS9StmRL2Lg+vDmsMZxvnOQVGemv0x
7dJToggGhX5rRY836Tt+1j1VJjtXmavGROteVbFyGcWpS1pVUxLwgTFYki3iGz6mQSigrWSmtvlZ
sLKqdANwZJmKH3jSDa9jkkImjyofBRszkYv0PpFld0IrelP81vHSRdWfsilJ596MYoZuZMEJJmE7
q+aidrHyHoFksurh0Nr+bXm4AVDYFuBVPJffMPDPfH1uqeyMlJmku04l/miivRVxFHQ7mVX1rAUy
Ue6Phm2AhmMUl7x+YwgIt5pxu0Sog/wU1Uj4mMDXXbCB3B7kD2CU2R4aXyQUUGoUS+648DbjtjMH
IqbO6SXyYHGVwspXVZuX3330fTCPgJUn6la9/UzSrzVhM3M2HeaxvRpjMVeokfQ7Ddo+ea0xN9We
cO4VSV7GX0bru8d9lO2JpHmDcqLcKjeDIuY5jXhOjJLP4xQQQmoPHbab8l7YZjwPf+xxZw0PRagq
7/7VpD85MNW6roFb1U+GpCtxdSbK0ssc4QLd1Ky8SNx9z/VvH3jDApSDmyRR1+fhzrP5s/waqE7G
pmAdeVNOYXFXX5UjDSkBynC9k3gcdqmVHjSkMtyztsNRkoU2pt+dTf0h3T4ExReVGdyrBzd6D62p
97WwZAvEFYHuCvW68kOO6dk8QOK2jzDSPrnmDVilM8Up2uBj33sKMIenGmE9uUus9jvBXq0RGag/
GmH4reOsQxVaWUqhe2tmvZNMRYfvp+5gp0H09j+Uba1exFippt0ogkaEsozIAUIwexoEbIcG7JM+
mLVWS671I0o4cPju2lhF/QMUrpE4m/U8cmJFkFlo1eYy6a3ZQBPjm1zHVparwY7318/YIuVTNbhC
4LG5GDn6oqmYYde0bqXOnZ5PbZKOu6mW8UpuWxan/cUt+q/yYnLx2EgcF5gJRQIS3dj4usNCKIe8
TwN1tr7K5QC4ACRD5CGlwWYN5h2AZqJPBYu6cFqVgh6P/DQ9hZvlo/fbP9Hr/SZukTb80oINZ9vB
zsMQ94IE6XY9pdDj3jBaNsHF7hms8mAFf6JdeLfmWNPnPKlWhk+Jk4NHHEA3e/iFw6Tb3GFdSegx
9xz90LA8wnEyMBw4X9zNRgd4aOQFpP957FZLNwvynnAZLMOmAxCyVrDVweOfFzeVvE8n+0jDx5nZ
HnJCc+Ckh7PSrRj+8RZ5SO8a+KBgebs2xLn2UTmsJbpxDYuHXDbzahH95mnXb08jXpw8LTpYc0LD
z+/GnRN0KxCDNlU7Y91hh94eMVQyivJuVj9VLrsJ4gbf5xfRe9M5WxyZ11aRhsiatfJFgSo8viJM
X7iFT1XnGAfkxYr/UCnBhGfSEIXKbSyzZZ9/aYXUwq+LJER0mnyfwIYbZ29UUzZcJEIlXyieu4Im
35tSGN6hS+VvXIZdq62Pp4MrMr7myFl6a8ScbNZxcAV//7QPeUkyCdgDRESi/BJJaWSXyn2SU8Pe
ZDj9CrJACIS8QRsGkw9PNBq/Fz44jSOhg2WmhzsCvEVughMmScpAp6lnXVf+Ghbp1weGqZvgxC4K
jZqOvMXjil1a324cHG+LaL0FOLcOnq8Ov6iy+38DYtgno2FWIa6Sdc+cncO09bztchzFmIo1Vqx+
OGj4jJQCWKdkehPUU4g7uT7Gc6uGi5xoPtPMzgFDA0l1DYUMjVsdDNctDRhkFH89Jv6w4r3abt1w
9SpPljjrjxwtE8nK9prsey9E8T+w0DnNvSGfAWHlLcymCckUZpsUojFY14h7mUkV8OT5IVAel5BS
q7rs8PFE1UQeuNamHk9mReDh8oGrX2DhcBloyuWrxPuOEM4+Ux7dcnrM2oEHJfI6CPyt4c6JGn3C
UCNrW3/Q3mocU0y8RLD+zgaiYWnthmrw8laWT0+wZ+4EO22R4Kb/PwZ5XxIKX2Uj79Eie6mePklT
sflGUKOMp6NBcRfZ7S/yZ6xuIYX3UB+rpXUNKBuAL2s1Rk0Snl7TudubHsGSkspCjoX1b7hMbV62
wwb9wBRX8/cjAYedQmU+ysPQjg2Wuz1J641AcAOveAS8ehFIstRSIbgJJ682xXSR+f+f7Z1BywzB
aTZHTccVz1+YaZjgBIIyFfr/Mjr9MgM6nOy/2KuGsBDBQm5hS0qLMeEAbl3JkA9+ta5nAMrqX7DD
FNHqOxseyS74X6HSfsh6vtV1bT1Se6Zz+6yCj40MccWOevnubjsVEYqxdSY1LLeY6AHBt84Rz2E3
UR71IAzpNpmGLCYvjy+aXLla6EbLMO7HIJL/3nOebynGt+8lsHbt1G/tJzlK7DvOEEQCIzPXBemP
MuSv3Wz0xHwovEA9PGfKJ2X9vrBeFHRyp/5I6d0l0rUE3gGwSoCpQilrxCKKj3bbtxcTwVYmiQyx
CwdmRuUsD96AO63mEuJQuCAPtSYRSNIpNMQz0GWZHagsrtwTi3m7outQzHSBdI/3VvyllVI5KqHJ
iRlE5A0FY7tqLFc63gUE6qnemvZb+SKQCqgoQBIYzHonqfP058yxm67MI6WRkXYXuIDY03eXsIoi
vf3eyh05TnXBP1r/I6yJGo3bmAUd9iWmKP3oWg4uUxW3h1PkwLVcrUEoDu015H1t7tu8Neah2XoC
s8GqD36TQ+pNGTjLronLs3e7WaZpPXIDPEUzMTEdWHtwpbl4AARFR7wp97pPGhU1IcMKJO9kYCbU
qGH2vtENuxQVN7xmf/7T9HPOLx/3GNFLWVgMlthpg/ihEiin4vGPwscY0eRs6fkdj2JRIQSVnP3D
IjgX8RLVNUKBm7+NBjSafaMRmQyE+7n1jjUeQP4NuaX5soiRjLcpd3q0FxIWPlQLSW+JTRp84LVT
3rk/JOmpdla/B6II/IUd9yQC4u0ZiWDfyt0bA6DXlRlKcKjHtIIvz/+1RjQFMJr5tE5kFB2pPlqi
Wt/5kA0wROx1vEdS5dsZTCIlYL/E+ze4YE2Iwnb/tdjKw6uqeWU2wGrA/rj+UkWtSlpPU1F2Nvrp
3eW96NlPyVp8mT8Ez+T+rD3iHrQfWWL4zBcgN37LHgTK3tWvn2QBu5MK9oCr9q1b9OxqC8OJ2Czl
s3GefLSuCeZUl6E8oi62AKNRGT1fxIae1IUar/gucc+0IoIFYmaj9CB2lD/g5S6FPKfH0RO+JeCx
w5chybhJ053bafMU1oH3zbA23XwcbIjodGACvdWNlU6EDwtC/9yJh4Aul/8v307V1sR0rIUDSLha
q9CWymxM1YfKXlRLGDVKv+VuQhPu7DK9gD8uzHC3dvF4oyyIApzD6PgBUTSYrsf81Zg7Tttm9gkt
3nvGIB+NaVoi8GerPC4e0iShZOk+N2dFJxujzVSBgMcstl9ih1cfE51JtTKSPSd/73p8WkLXqJT0
lVL5xX4Y8biO8gPNoeOIFaSXKNhRiUVGgnNcXz5JXXgXdskAo6NLkM8j1X365odbvI89Hx4fHJt/
w+sQS92WAbc2tTbdfcQDkp+T0wKaWBaiz+VnFTbmuSr1CM0WrGBHfjFRm15OLc4jYySZ+oyyloOY
RLlN1QAZZFT4rB3zSaSmOmlg62j/QQ+VfadZVPqSzBmVemUSeKRbNdJYeb8KuLsZTRpkfXu9zvUL
LhU76kCsmONDsHAmipTHZliV4vtJp96yw4xsx6Z5+L7tZUIeACRbRVWujIy+emNvmvmbgzBh0zFA
R7XMJqMCe8hf+AL1T+6zZWMGXUiQ5i2CKQQPnBbJ/LEBFH+UL7MERvTrjdHMPivr99t9ba1U3bAQ
HvXkeMZ7oReTO2v6sqiuhG5Ff2NBB34EgOHK4HNef46LjFf+F5OVYEjMhk7nDCHEpkAkLhyPuOio
P1fxKrRcS3u0jQrJvg82gytjdtgUzU0Ofv6FpH5hGqru/WmCQb3zR/5n3nyEQeaErYez0VIfeRcK
ayTCAa3s5mz0e2HRxoGLNd+6xLjnn6GlkBqVETlikhjKIetda3Wn0mkRURQtub301laCpPZ2m1r5
DfOaZM4y8IoM0lOE+NwH+Ti1YdBbBBb1HIx5sKq7MaVWB9qEmSTIcr35aaPZij5eqd3SDaYr042f
HxakoqZq7XCu+yoGnmANQ9kjiqNaeVXOI4TYaxz0u77UheIcBDJmx8LIi32mgwCR3Ca9qJyVDVBM
V/GBwpph24/wvd1vdkF3eVLYS3pCRy9eNqqGAQhKAd3KiIfOkV+g3brMnZyMLFB3Z/M22iEd4jkj
QSmdqBgTUfUux8EtJz8lVGkc/Z1nwx0vsi7nTolf6SnOjZGwZoqRuP/yPMe7uQtGGn8PCFaCQuAJ
9a9yOFgErRyuosdAVQEm46PoSBMpjHZN1UxD+Nn61DaT8XxD/JPjdc/p8GtayosgXGuM05WUKVz0
QoBcMM6GBHoYmrhIi/o4rgbdWZ56/u4CWMT+UNbPX7uuRa6yJrjeV5j+2KsizeaN53DT8WdCQHyB
UlvAMxpZpYy+B+HxnQuwOXhlQXplrI4/K80htntd6WB99HY6Gf6/Bv/GfcbUA0I8AHji8phGHmGh
fUiPwFfXDJPSs6ZLZY30VYBSlhOFuTzxaQi7BEBxrWy1HBBP50LUmZhOI0e2MCaNUic/T23GZRXp
QmksvjO5cAisrjNQ8Vvvl6VzVj7UpmQNg0FU6tLmUdaq7swYu+TDr4tRGOx27D+4mdYBD9IJBxK+
v0gO0WoHvQC+MlWnq6Ld1ziNDVQ4HG/jUp0s9bW+VUZEBkM8yfN9oiCR39ECO2lG7tEiL4sT9sqW
SN5xuvIQEENQCCBELevxWD6qR2VMPHsFsagG8zSH2cHah0qNXXOtdCSjFvMxY7TBqE1L7sa94ElS
BZ0LY6QZtizGvpItwcg0vv2Zg91bYslzVJocRoBdMJzzfbw9JZV1ztEMbmRu+mNthMHQyBGpu6Nw
+2icAngl8Z64y2dROl77jWiludaqj5ttGXFJWE6vRY0NkiMfvf2rpR01A9X/g7nkCnmeysZfKQvY
To6vF/CYHEqA7GAzOa8A4pjttVB289BL0GYaYSOPKS9tJl7VDo8Ra1LWQ+q22s1MAo7R2hOFrSQ0
Urxi67a/n65F2rR1zKvYBS6YZ4E5gOqOnNGmUtcceccvh49nwzHqe7HS3N/cm/zvClDVro1fe0Uk
872yVLvfFAOS15nTyDKj+pVCqpSj/s37kYFZXPUmV8bdh4fOjd1Y/RchlxScr/POKhz69v+UzGKy
x+QsA0kSUAtRQlf4i/FVcRXJCH0QQ5/I1E8ifeZ5573gjNjdMwFySXJp0jjtBdJOdEaYnAMoNr2c
naxqduVfDU+I2mT6QRxTF4PHPN+yr/cALI9t3LeYLJ2tqjQofr6QVbb/1RB5rkq/DGuRBsMj/iPq
NE/sErmrT1eUtpyB/jTVwHf2NvD5i/fQDadOYyeQSsnzZg5iu73EPW6UJxnleTLxu/EwtCOV8nU3
BudtDLc9DdOKg9nzKIns5Rv0CV/AX+Qmj/MgRzk2OUXvBYYXDaQ/K9WsgFNV85ddqQ51SmYix1MI
4tOAR99/bB5KH66KIRfA2AqzaZjCgn8KbgzrH+zjS+GzFx2ee8IK1I0qO4VwjvD/DsXfNNpiTvvY
inigMkuIO28C2MnOCRp1D/i4Bjd4R4cAJYrtipvUvdF1tBf3eYVkJliq0mPJ9Kj6RN341/q2WYIP
7Qbf8SX6qeofYFrPifTa1fuz/0t3/75xY4rUJ00AqhYD2sXLWLCEUtj9/j1tiMMV+jmovjYZx7jr
8jfwjSP2docOC70k1qLVN+sacwkgYwqKrWhYhIK0Y7FXBOYhjwhdD7z8kgLNHFS+D3+3prqi83y/
9UZuNhP00HwV7ka7+Jg5E1pdMTBD+P2ySx1h6RUNF06kKXYsUZbTiB0NKd92KhhPsTAkB8lZMZRJ
kOYzPujbGIDb00bAfn8GN/BWgSlPVxDraGCgO3bZhydR85jXSzf8TtMyMpYW5M+fWGgDxyi7fqCH
iY7UjpJt8k8tqKodxOHSiU6vQIVoU969i0oWHpuNBriZ9nUmysmNHwQyravaX8VG5TLjXyJolfFk
EApETVtnMtENgBT3FUWdZis2Z0X8bqAeL8wMv0eoWXTmJCkfHBru4bztTxQ8kRbtsMqWcS8sl8Gi
44I9l9sYrxhe8BFr9GyTl8NQKTvfynSo/ayfGKXWOF49THjYUHAHiuA9ICZVtyPNyWrnKzZAlblQ
CpL4UFu4Citwhid2z5tH7TXHIsoL4HidBa+c+KYqgQ6b0GoEEmwVMnATWfQ5vrFnLA0XsLLtSHxc
WZKmTKE7DT2LTHxYBG752zhOZ4zuqTzJQEcDM3Sq44DG2aSCEnTaMWj3tqNnfsPkSoOgYnki4EUd
Z/GTX1yvw1PUPNtyIWcd4sGkk+Myk3lhkSRA9KqMGmr67XYS2NySchrQJu44mkGdwHinwEcHMt8R
AKFF1fejHRNz8jbKEQyBw+drzmZ+e9767hJ9zjorI2fpvBzOrxaxMyJOdHM7R0PN1jKRhVaoa7+d
4lavqc9qEnzk9OXD3ST3xAR+QOY4ge5PHxv3EptbG9/2fgpHsqdgK3YZCjCQR+++DLyD1JvuMD2e
UxH+IdABUSh+fzNGf3mb6wIULQP7p5U0S4t9GxdWpjEZysIE9+F5/jI5mw83Se8Mi+3OZWePWl0v
4NGcgmS0GTn6N8/ZVt5qHsg7eyij+8x+/v1bZu/qhIcss4FH89k3oPmakjdiGychoyiyL+CcZiD7
fqI1STTvCR7YTWQBGI6euiCVP9qqDmAHA3sWXzlyucKV2/LVfLJIdiCa2YE132LYE/Iz2z29lyu1
nP3SehNuSt1XWm2OW98CCf8KdKIe4ag74A963TKNV0lovFqnXNDhgzOGh/NU0Nd0HHBh/vb9kObx
/Ddvngl9W3LnvQLWozhbWCak3RNi/ijPzrXfxTMhNkrtmd71J3axduKYCcqECiTpvcUF4cafFV+P
a85gjASYikYygKuw1ISuzh+THPnMIl17dprFfQiTr7uDwjcDtI88etGSWwmD6JHpamNKQXfw2dwB
rFDz6QKVtQ7NuhkckcXzRhaSgzOqg9mOkdylzuTBQUGB4eFU6u1UB5vsj8gtGifT4PmT5bkaxI1B
afwstPfe/faWUOciwXRAqffp1ANsndmY1RRDCywwxDe/lftN0KYBLI3gOqNQMhQyPdDBs68/Iq1A
l3s/K/Ln5fTL/9ElK6gZLDuUPG5T6TE3hX7eq77+2kXswuBA512kVomQmkeGraFWogPExz0KDJxC
XGA6kbPEu71bqAAU8O6BHUDu8OR38aZhnEE1usRzJf/Q/Y33KGhODpwawOWrdoNS2CxBnGD/VYCs
sCfyZ1Hi0loiuduE2qWbvELwX/dC6s4AH/c7cLPDULZKXCGOliIfdPZlTsurGpIlQeIgkhUPbzRe
04583p6WLcV0yhE5wLZeFph5QswWlyTmo3rqzCG0dH74kXJqTHYB9CD1FBlXsDKuIeKKn91l6slI
RqfSWVReY0+tcJNTx0AAAHas1rccKMOFjJeEUNfS7Fj5Sr7QIoo44SogT3tsZHxTFaCHt71ojaza
XjVhvs2forVpMFhdbQ1mZfTH/AqJveEAWs8uJaN40T0SuJqFbhJy63N2tI0TqTeI0Fkh2bdnhAD8
4t5SBaXb6EVghbHSHLJBYt6K3amcInuO5YSNg5SqzzWVFaK/j/xziRQdeqfwWHqRz2bKfUlhXC8K
Gts0EYUx8+NxTaEV/7cB6OSb9jqvFKU42Bv2NTPo9trFTaG8pypjlaHIRq+dB9ckJqhJvlCGCig/
Z0cxT8xScM6yPjjhw05wk19HJyZoCpAYJYcnk/HmL/4gW3HoVpbMuX9tKTfY79PMmZFpTr+fNgJN
mySktwauP3h3CN5RurwETFsy7rBPMEQQsDOUseTANHSuH4wJJcJxbLve9NF1u2CKuWbfSvrmXarC
iWdnvjEKWmph2UBS3XzZDozi1pryz9HTxOBBEBt0xkI47HuCLSj4CzDiFjNfSzEHvWM3Vbz28hvm
9St/H+1ylrxr5TZtpHsKKEc5/OGseJ0DDJ7T1vOvZ865bCdbB7u1NS7/BHsrpiyx5hvj6qabAnHp
kdTiXWyQBw5X554zU1ZGLpeJ+Ebir1sHoclDygUgZ1gQ93FgqwMGJm+Lqnj/GHgfqvn8eGA+b472
4o9sse3ttuGCOWS5GsUT9+0btJqIjLJusHKsNXMiX89XkVVK+uTqrD/jZXyNU2wXvC+GEhYxoJ44
S0r7LbGxTBrv+ZpLKrkZFUDAPVXWF1PrDH/VT7v2tHhnL9boLnkLdKK172OEiRq7kYwC7ocuuTkg
q3TcoENXVOTuExhqOUiUl5/52Dpxu8Nw1jIoL87S6Thg0zK9gpsnJrkmqqtXV9VBPCo9ncYtV909
L4ucTI8M5Id6a6HNs1bM4erowpLbKYoAHzpWgcfme4mYmoZnJaK4rAPTK2gRpUTpin3Gxxar6xIx
jyPttWUuhWZD+Z9ENnQKbz684DsCwXBMBMwn+2FIe+AqpMgecYpdnGhPsWZfxdK3RjKEAEbKmmQD
q8Fp6ZL+QPZyY5qnXGvKscStaK8/I5fMfoWQwIhOFRkQf5N6OmP0SOKKsH4kqNLmdnBNxt5frBm3
sQ9HSZXXHCyn1yRPz7jHIQQxS6awihILMM0JsXOr244PIwrK8JWGoum1UUTgHZujBuet/0jAFHOv
UK2IVoJI7b7UV8mPavV1mUxRxz4E34NFK26bx2gPfbgCDgqjmkDovMOIXrScX4nRhjWk9jQm9SlX
SPKIg9zfaWOc6Wh7FnkG6DfLv5pj2hL46OmYgWfQf/5mp1yueHtkLTzx8A33WNWf5zf6ynQVcTRJ
N0XhDhmOxbW4VxquKaQEAl6BeX72poIyvtZr2TXIzgg7+5UNTbc+lGINmO8hIaiCXjhrSOyyyWp1
Rw+ARLgHhdvybQUInPXnmvk6Z8f1/f+bVSQVyAtGMPZefGEV73PIHCGlI0MSBf93+L+tWaZvRuBm
GDWcKYg5oK9bIy18oDPP0B6+oAzME1N5P7opx/S/iALZtTJ1ooj3oFy4XB4Y9HFD91HKPHTpnVBG
oEbengqrXFSqdGHuWCtOmhZweni5Fp0P2GWtonv0AOSF2Q/2HRd4tSO9BpUkke5L9BFngSLQA3G1
fdDL+ge/FfsrUwlcGlD1Xefm7KEv4WrfpbAjxHJ53d2/L0cd1frd63AH2Uh+Z/gFkHUfFaeehYFt
ngxE+LKT0dxDhtwhnRjoJJwpbeF4Tq/HJ2IW+nEK90o7dsWr7mlQorBR5XBhrYiBcPsBZz9L8Xn7
6RqIFlyb2C3AauTbDOsHVQkc4l7w4WncWIyWP4AyLuUen9fsSYsTVZs9SO/ratqwmmolDhwLNVvQ
51cVle/iaa7OFWPzxeLkF/1EyFHj36fTnN9V/tTb8QRhEszkFNuyFVHob+ZqSp0Bw2JhQXRgBPwq
5u5KWlaXo4SQ1sVdmBNthtsYn+IxbbM8nbaBjirtUyE0YBXCfDXNIiKStikzgX8A0HiSm2Ap0YSJ
nZ6093liBHwgYci+eDpznrTrQA4RZXhcDUMtkUnXI0m/y9EEt37NkYAx+q90Sio6VMBPGVnFMZOx
yQxO6zFdkUlxte5hoZfAewZK9ZulGLRRf6ntJQ8xnqMdbWqrqFul2xQY+74phaRCibTKHpt+Cufw
xo0XMmf+K2WLMdyEEocm4R/kHEdhIgGTYoi0LGGm+rIW4C9lO8KmUeWuuirmh0gbWXlgPELAu+Yd
pzgBEpiMs+r3mvxHWKkH/eVXXTAwO4fj5ZPsf8Xsq2GXvNahLHkeku4pevRLVw0k3Lhu9riS7DXB
3iZ+sEDZJAR8cBnfWxE0t2RQS3icaWgAbI35+ogG+NmCSyX/ygkX6CzmZcgjjaN2lwTz2wzJhEgM
BF3HBsUB5ODcrr7E03iENxrBDSIUWDtbGEf5FZHVWjnVvCQDiS2nVXHjThWM3c98IC7MPPabet9e
eecSTAlWkIAmGB8enoyAXY3s5EKlnrs69UuB/sfSJkIDq4IG/XhxPyW8aBDlgkc+TxxuAaiwtjrS
WY3ZOgx3suh3aJ+qvrcOMOPaFNkca7tMap/POyoK5DI4SOdlIxgFCoWyaOnxwgLHjq0f1YwfCJJp
JQmusdeKff+EwKIoo+KXlVNFnxqspjK9CM1+xtuuf1IF/J9sarRKjRIRVlJ84eRNagOvF5pC/x06
IT0QJ6l+Ff8Dywwdh0sWhcXQSt78PRCcnOYIdWpd5kVYnpcrofhZLGiAqlIszmdTRjMx9oAltCrV
1qZ/qkzWKX1Uu6SsbZIwHzd26c4o/JoUpQRmLRKxAUNSHtPPnLTQGALhYPJNGFdLjJI6PWqkYw91
J8doUA3iYUO//rSYwywALWaQPmNE9zcjkB93DWO3fAg8+LzkYN9Lv6dvQhJ4r2m1U3pFDbt0PKme
DJSlsTx+wNT81HOAGp/aCC1Pmax7UZs0LytDdI/VRgDwCWgMORYd4OZefh4NwIteWf4TYE/82ppD
4qIeittuKsLGJuefgnjFOgjSQuoEk8LB+ithpHAMRYQqoqLT7VRorXVdaP/37elfIkvtNaI81B6N
SvT61/ISVYCX+MtE7jqdCxv1b2f7gDZ2whIIsVSpHQWLbfNmYRxQHkdkX9F9g+bH5J6DNH1mbW/p
RuTZf4dwQOyAHruGp+IzsT4HOCg6ihC7wvkGrBqJtxljQ66duZ/8L0PtIC7rj1b2Mlv8nANxCyF1
VnNhdrG/twF15ViNf1c5UkpOEtThC3/f5XMc20BeD2/HScj/UMipBFEDAPeeHSaBduiWIZM0O1VR
XXciAk2c1JjNg6SKJv7fPScPQPyWx9BFSq0mjdCeZaE1pCay1XEyE/F0E8nVhr7s3vTlFue+9sSG
IWnq1mVzf4+4L60v18YnBOy/yeUQFllGXZT0fY2WXwuTsq1C+DUoW8Rs2aspMCCk+n3FqPrXs+K4
gZnLvH2kVjzl5h95sxGe/qrD+0yAE0zhWaFYhuINJ9YXk7gTLdrW2nuBU62606vlPgh/8Xs8lE/d
aPIDtFF23WltE0dbWZnpMzkwSzccZbsxdZ7rJXfzNFtE+eEG/R2BoSM0lR6pD7vmKgcrvlABY50+
Y00R23tWkcLkzA2ezOtRZqEI4GP4XfYChHgsg1VaTwslmAt9xjSh6DwvrLfqnHqf6MEopBizVSwG
pnt7Ah85RyXiQgz7lgqcMVQOfeidqOMQcWPJolyRX2L2Z4lgRqOeL8VdhcCbeW3hsjx0p82s5jxn
qPDc6rduEWYkYaGh+Ei5Dy6tbdZzoCp+gVGDcKGVymJCU+M132+fKFvODBRITqwvJ3VwEMF5yqmo
2xGHoZq/pSiTsRFl8ezU4ArdB3tj4pN3P0AG1CX21F8v3ubY5Gz+X4+NpH2yydJoTaCFaYOMHLeP
OT5QnTvhg7RXPYOneI7fYGYA7ZrBlJGQAnwZPdoOe+D3Prfy0L7YZrgXc9sdxPLVejLFX8X8v/Ns
MPJsjF3/KgDiEVDG6vOPnexZjWYLPYNr1p5VBL8WnqiCkI7uWqtArXJKC34Y2R7+piSi98ozY5gq
FNYUikDTgDcgqqI4HQVXVHV1Z6j+4MiDDvGRC8YeRJOo8sybvk0TirnfAtpNtEEQVewxfcK9zhfs
sMb/waehLsDRx+wyx14cjJP2delVmnWtMLmgJ0LCEgEyDR56SNxT3wsa8p0u96WVG7unh6W3jDzY
iO8SOlTxnK2XTuQUGcU8INv3iyGfTox30r/+25jQ6GWjFRFhjCiTMvJPFDQ0O2Lv7LLv01OwXx/B
11ddraWysTkB5PxpJknn29dHGSDg3kCY9UHnTGp0HLaveMHwQ1Vvk8bHkJ4lL3khIrh7yUpqj6Xi
9f3daNiqU1VE5u4jbkEqDMG+YPcWssTHZlU3RsbIIuhPbNPr/jReTHLdPtS8lcDmgYmvKSccwq65
EUqfQ5BEI9H2BAuLsRTg4yukpEX3wWP0DKtIWp77uEi3wu9tYsui2G+UxCMxRuWRPmbl64n1h8Vk
JSRcslibKIW5Bb694KdFsPqWg1fny+llV9Zs9NYvfR6Fx2U5cauWuwMZk4ThgJSEPpJAxoweNm/c
YWzfiXbEA/TpAnne0VOdLDxoB+MiHdyHgJOOoE4z2macPmzW20b44RHj4CaT33Nk7bE620SBPIZR
v5n9m8lJ98Rlqt4KZMvE5RyGZJ6LcmAazq0GwBkbNGCvZiA98T2uB+58JvW+GAsZHlucq4oWlmAg
PkgCaYENYorPXRykja0xruz+BBSgAtzewJO8RUjJDOTZo2sm03g5EZUe/khdtqEGoqco0zSr0JCR
MZi2z/hovngvkRXi+kXQI5i/OktSfN8AX9kXqeYp9maE2Jxo/KILjipwG9/UGps65Mo2FMIjnLX8
DoobZzRECFcc0D4t6dXpzE3bq1Ea2RNlSexvAo2Prj4gVUBo6xlpc61HW+AHyFm7PYSn5KWHIJLQ
ooOJDLvsHzMdMVE9f48qh2H6vykNwHIb3RlhDnImhHfuXDrBkiuk/jhKLx1fGXbAnMAE7/LcoEAc
zGnLBdsrROkBfgoOVlZ0gOzzkJ16lEPep/IchXb24QVvObXhZziQyB5Ouq2i0w9fOQvoEDU7ocCw
1U5l7aeD5SEPIZuq6PK2yLP72oY8iqKnJB4V5xGs+YeM3UREKuK9CJYvVIQpsFvtvgKbE+oRY+/H
jLdH+beUFQaeWcAFwHQyafa8pyBq0JaVyhAB2/XPw9zif91n6SABY8sh60cwqptToPNyo9UbBLMU
OIF2HDCgPisFJ6HYXQY1y8ZPvibvPWPphLx7rMbG1CoqEp8uQ8VmAnosE8sJxMJnzL45TnEJlT05
5KG7ZSAyCQtjRgMZLezx+LQ7AEMbdDbf74UH5xyPRXqpf8uiw0uzkTl6lW/EIehDa8lfRjS8klCe
pMT4FJsElw+WzNoWy78qD64vFu6DOfJ2REsESyS4KdwpjipQ9KFEiRu21FlrLWCW7DmLLtjMgCnl
+szqgW5UaKW9zAM9f6/H414wGpR0O40CYg7+MTPh0Km5H1YKbcOqQXx1WXFmOjidnooJwT9kAvkO
tTOmSXd+QzI8o8w3wStqKYxP76D4y2fsEAWYLE7LUNeNhG9lJuoOYE7kd0cGSlBUdGzdkRQs+exq
WP/0IkRuwM6FowgPWqP6aSXTyxDun6GU460mHizUaDBkEfzRBzj4UKIXIsxO1f0MnVlSiMnV/kOr
MuEH8c57eD7bzkvbrXx00mDcDt/lysG9vPvUFUbLNV+3Sxy08cXzkiA/LV06qY3BWphbcQXmmYUo
6SbmzyZ903KDoeeUiF1Y38llRuv6uMNhJQm1IYVcbhg8r0bJSa7acE7AX72W565RuenqnVSYFtyP
NEVIDMLT8ek4ZLlHGV5HgLYjHg+bfhEhMXpPR7bXtkjl96YLAyL4N7uDUiCCQVCqIHSpno7vgjnT
xmsLnFtzJZLjIwy5jnKsg/o3k065aAbTBkBcsnL4C+KnykRhVsmEkkJYB3PFnauhbCuONCF0UEEC
sO0RhjHVbF79JewVbB30Pp3r97LpbvBVOylURJh3u40CDZUmJUo+/awzBXrLWd+qB6Lo2oOQ9WPT
TwNU7BVr+MyALsmW35M3GH5a0m0+Xv3K4cxsJfbGBANa/E3DDhpKsFvcnaU5gfZtnTFNCP5V3kUT
o/8LG10X/Xt7qEP/4qS8R+3wTqGgx9tA4CbSNEJKZLOn+KQs+vge1UBcxHdlObbdTNOxWQt7fiOv
pJcjy2IT+FLG6offxwBAg0cfmFhga1HxncLidiuWo84LVgJDiQ91plWCBgaBXJ9yU+s1jbqL3tgZ
qKo+bfKu12sYoLK5h0S13CDX4kWIdR1mMkPCL1FJ3MjVX0jv2LXtfeCV0+2tQzrVpE4OGolZp7Qp
45v+5nJBKLvqv0z5gOBiem/y/yxLyDMVp8Ue8Vxga3qttYogMK6cD7WW1eROhEy34Ty/gpxIbFg+
Qed46HDnU+c/78csr1XwARoqvfsCz5wcz9mWlM5NxAbUrjSPIOikqLkOPgJtKGpV0JpccmmfLT3/
J2rbDQlkX3GMtF6BiMULWqMqc7LeHte1+3VZp+8u4g8iiEmOUYucSb9714+j+bvOX1zf3sd104bB
O29Z/Bh3OqlxQdLl1VFCgSwT6ZhLrUyEfPOOZgogi+C85udgXvnAUsbV2ObhkpwGglDJCvlVWT42
XHfm5Adi/AgB4yMSUrGuIfTSmkou8RQ2OihnKv9rr7zf1+eg/pKtrAyD5X+Aks1PWePdnJKfQAVT
FJ3xrXdaPw9O05SIo0Bpi1496e3rarC90fugoVoWpMfxQ+4kOqTVW7dO/Ekh9TTquMjPaZCLzjOW
RmC8lf0SunRfJzZsutzQXFeefdh/BEm0y0ZgxxmK6qNKX6lWiHaJQ9G9YD0yzhXbz0ej2xT0vhCE
46H5IL9fAVi0v29XW8wcZ5JMvUeNfICgyIhTgHitjxV2YlbPC+YECO/q+17o9KHMtEZf4him35+y
7qT6coyvbyVeB21phxnAAJR5aZEC5O25Xj1kKXAq4rGFhm5Wa1gdtuEoI7kjBBH3Ajy079yz2vAJ
jUE/WnZW7J1rI8ryRLLKBfPtjvXaD4LUVj73gBlwy24ZxSVTmw9kwMGaGREfGqSnLk8jICd+jyL0
nworFdxBxglbzWIWhC7gGR4mkGISPkQ+zNVBKxJ+DFMVgr+LLvv4aGcqRiNOuf1+AJzDSpmiBMhU
8NIGPCvxnnXYO3YwkRd3udWdQbnOqWQD6mfyomhqRvcBnPFj7kz+6aOpEaQiGDaj2pGEQ2aIj2af
nZ+Q7HDMpO5i6I/94MKTz2AUUT9ODMHdV69wUTr7wttH/x4hgVVYD9DEykTaZWb3E4uxEOZiSoyA
Im/48X3DisksW6vGV77z2sRj845TmCnGFsGkflPcmrLHsDF6eF/MgWdZSx2UcTmjJFNyKfG2/8Iu
ww3VvhX1FFKWjAHEGVVNCwqpuwk2IacpR6XRXe68nzldKxGaNCWr2e452TMXHqeHgKsLauVn3sRS
3kWWHqNCaO95witd6BXiisyflMHKxIgaL64bMzY/kktIw/sdXNdpJTrweg6BqGxvGsu2Wkhmuet/
9OlrRu/2ah3gAwL2Hljg3iCOwuP2/1iHhXYAb0avDuBRnnD9ehy5XjQKQARHQMj6T1neCr5TTZ3a
soN7i6soHC22lyiNf3XIOKVkgV05RhHsnuLmbwwqz0C3aiQo4vP/GDJN04WT4jzbKZM8ijJXiw8w
aU+Xo8457H2mA0D3m4SwVN/75r+GyMLsZyVOqLdvz3i5Z0ffLV6HLLFGX5nbuELuwDeg/zMq32JK
R2oAHUioNhwqIfD1qOvwxHivhldj0DSBM2nXc0Oiub28a5GAcB86JbHFl8m+MY4Y8Hb8ueHV0SpQ
fVh++eCNoStwI5LlL4LCdmODRzcsti53EvBBh0xMP5Kk2UWP2yrFCy5jvibEle1KRMYZ8i5jUlmF
uup7K6e82DhjxXj3ewRNXIZQ4DM7qjbBSbpz4PKBJt7HLVYu5uLCm2QC68PlFzD8lTEw4zeNdtQT
1SlN5dH6uG4C9UIgI2V2lL16EgWD/ZujpXn6ZtbFVJdd5weC92y0cyixUpvVP2/SJLzikwxrOcu6
/UrxHI8kF3McxMAdWm7vSCARADsYJ4mD9cFP/q1KHebMtirq00jRDU8VTZDCoKMYZV13smY03u92
MkUd4fCr6UpBhLsc2KD8zvSJykUQWMcroPDsxwduufXO8s0dbYpkCqpnLwJeMFCXTutuuKzoUr85
xJXHK6qdbPnycNaTHx5IZI3bDH5/LoJTluvBAM4+QypPm2hbKT0yMxZT+nEaMJn1ssVbz+7lbd1L
M/iC5q0ETq5F0q2rht8FAdTnqawhoEao1Yl5dT0bkpdVLVwSCU/WdnvXU2WF7TTYWHWbTkLalSFP
MesB1Zn0OWuPdVQJi6r4xEYpJ8gzWdL2h2KwZGNpO5vyqwlmZ5rWh0YoyMOAZgNApmyn+gho6TWG
zHvQYUet3rrVLri6SaTusjjqCQBK6M1csz3qL/zz1fzplODyBI2T/UJFn2v4Enz+rCecASf3lETW
HWdt7FAm1DN59gAw6r1L2YfxF4WXZnIY/9W3I9zMXKM07iweo2qkPYuny59UBOGGc/8WTqATdqkq
GWu5/0bJQHRIfZcS4PYjwMxcrJ/1hprg7hIWcPc9n657/DfClwfcZ1P1RTvkZGU+RvyKayGOkYTA
vL/AesQ7+qORAa7r/vHXcdO97cJNbbkSwRAa5unInCBTtEalfZGgDUtdkbHF8JHwIIY4mWTPui1A
t9faDXcbSBY23MdYb3StfgyPM9FIFs4O5GhElGWxHCRI29n9AdWn3vVWkDbLvW6rRmr2tLZEluaS
8Gw24L8CX9zuw5ydWv+vIxPyP7tnlkMqfN+saEfsCxzd2EPmrWOz08wqwZPj0dmmq+uNKt3EbZiy
CTiAGo5UDgJ2Rv+CrZz70VcairpIW3oTPFuaR6f9BRMD2NCiBbyIPLOgDsxFb+48oij41K91NUdV
nPG/lAFh6sH1ysM9Jpo9dzZJWhTP6LEbij7uhXwPds9JF3BC7ICuf5a265lmXwfLuxVOczv3ZC8J
qKRL/GOgU3foDQ43VN69HDL2ui6YFVGpenOJ57tGA+ti3oyRGn3n6qknqCRzQOz7xiPKJDYTrR/A
a3bhVnLqkzR8JKuKitfZTfbQFiqBEO5oB1RArbssWAQ/9L372EYS67Pzjn5v3czoOLpb3ymoIu35
zhTQUkz+TbRB8AptwyfONDEwJ42nZgxGMwTQwnx5A6ax+O4LObjSoR9PYgY+kfi42cgwMhUK0N+K
iSE8jWAzdeWBeumJ7dYnM6PUaObVrOwXx5WM7AtyuLrd78vKYB5RAGSZxlIMaNn47uQRJFMvr62C
XQRM/IbDfiqLJzz7qlsB5pUf/7bZoEw4U8rStNkdK+4AvEDc59m51Giywaw3srSr/3P+a0xpcFre
ZCFC6PKGjpQvF2o4fnHfrNJ0A18qUhILSB3DrrNw99depDpCxfH2DMcAzDnpVvUg1xx8/fmyTFjH
sUZoQuDOnts60YMPbXWw8s1mcXtevlgoYJ54xcxOeun4XfnHPVNNjb3nvlsbY8PDqAYaNzDxAHiq
YdoxPjn+sX8l0aFpy8uhIjFvERlhb/8D5n4fC2Aw7AAw5GwHnaLCPjdxFGkigH1mV4dGjIMsfD5U
PjbbS3bAy7DjdrmtM+bx+7G1nRGAHVw/DXZOA7zjjbBd8Vjbm4zuUBtunbM1x5vZYr05mBK/Grkx
LTsdip0xQ+JQZ7Ny84ycvUirU7UAMxifB4QZ6bvqeuO/ijG5JAEkzAI+9mRed2hmD+5RIBLA5M32
IEaz5kQFJRNXCmkt6Tg5vEaVOVwRMUsnnwztfZSKjlWCg9N6RU5kYmOKG4DNDTcfMrpJTmyFgr1l
oh86VDmc7/4m68zBwBQSahC2s6EHj0eMs9R5XXc4WVkayLExMkm0Uj5POyLqYfDu6LtCU4WObnn+
kaO6X7nQ9EylyILW/2kl0MtJUP7Mp/Z2qqgCNEi/qjdvJy29RLc2VuI6K4z0AEeCw/qOLt3F0Jim
RnsD/YyI63rFAS3heJ0tbIuTrURcw2VuQmswYQ9aa++kbpyef3hyqroXk7dCHzL8gBDc+PW5/lHl
xV6fLnUiBa8yr5BDr3/M8J97JOsD3e66Digp1qtyTmEhyIsKIHByxLFztrupsPtq+uDoEH/WTKem
1duVnrtUpdWSkPlCzejuDOdbGM9fuXbU5efKWYHXri/WoyB/2ND2g1CY5DRmMjMZtZTl4aTCS2YC
4Xp2e6WGBratjAVvfV4NwbYTwBUbzdz+idpSnRkSY6jYZZE9rREy1GxSYr8vTa54qbJW/D//E4VV
6cQ+u0pMYvARhlTyn4U9OwPdt2X/dFlpcwh/GZkkIXyJhgRVbEpqh8uyGBg+DapbC1hNBaMwJy3h
suU26NgQjgOW0+FfIP3Vec3AQZZR4+UmXsZPnggKvjdAuRf5L+05v1XI4atkOqrIgyfPXQ3zMjCi
m6jvJckI1P9E5sTbkvIdtUF+q2HYtnNGIBDDyRR9rqHD2XcfTuhfRPcWrFORyaBqUkyKqoytnTNT
+MiqeplDwNwQRw/3Jx7vxqc7pfgrsxIfhnfTKzejBg2vN6pmjoLaWEKtNBpJu4P5LOvYUWOQk4a0
ITZKOpcD4ZjXmwNseX2j6epkhni9K6+nDzLL5ps/3pyDH9ejEvsyw665fK1q+mOxwSLH9anJOeMT
muG5OJgP1o5d4jmZKLr1VLf/dBNfVX/ADECM9sRB3jSxOrHamcqdnAznrQ9vk96ZijHRo5nU2uH+
xFt7CH6Zl1JvvKCqHMwFNA9OM1d/BTjpTMVeif+hU3GM6BNGjmTJ1PZRkxE3iB51bh8F/+fMRIt/
zHp+sU84KqxjP8LF/wSzXBZvbwvaH4TbhDEnm6aW6XUnYtwYU9FUeXDWJZfTRk1evuIJVzX9dC1b
424Z1TrG2Op+YDAAS5DBfLISyoumCPqVhfYvAEtQ4uklhFasRiuBR5w9r5vghvO12op4RVsmqc9D
6kSG+XmjFm4M7xRnYFcoqyCQm36fQ0sYz3/BUWHy+4/qbpmHBdlqrcFGugUZsC9LYBG5FqnGaES0
GSGvbac6zULU7RZrGhiReQYjdnEJdtYRfwUFl8tlrN8+by0ftkaeSrC2rw86Olm8fUDh1738Lvxt
7vXMuS9GevC3Tq3AWZqYbzhTF3+9aXvxzqJzuTB8b+WzuxvtL6gP1EJlpimBsfpYWNxWYj5D3LxI
WBeXP9C9yUzrsn3FmhU8ojWi4t+VUPAi5r3yj6U3iowQFy17/YSwGJIGDr2FtIWzJW95SIka4+A7
kwMfDSjlYLdrU3nOMOAPzqYZ+W5YPR0TbhtpY66IiXTFfUzbVCNPZneRPRv/pIsjGwO5nncpyQeH
E8tOUOhMSenIFgS9aYROBTAZYVQIMrh2+1iPQZrBMaYp8ppNU+cEGwvIRO9ksQkDhgrUR9uWkVkT
4C9RzFAmYZnOAREh/8SSQAFzyuEiKHLOxozav7QMUjHWXUlCTjBadqyf/xnd4ySEnKQ7E5aRJ3UH
Ixz8gstjgyj6ck66vl2MRxsttXn2+IPWnHJiSziKfwolj2wc/Qm5WKZmTYF7TGKiWsU74rLtNZOx
m7/Ihu7dwzwjoNhdqMBcPW06OA7JivpuuiS3Gpgkqz/sJUHaliBUJahefMgWSQbz9dloQ1Ab9Mx+
lDzaG0mM2ww6snoVzSJXPbZzS0tbQnmjuvmaP6SVcRewjCr5g7yadY+alsHqadOmzHMh69eIdTj0
LsDt/uXPTSSsovo60ra93EjRI7Y42DVM3Wul+TRY+Afh3uFtjE7jjnyY20DnFFfIyUNazCEw/PpU
+pLwzAFUYN+Or54w8pwRHY51An7TfAh/elZwauyAM4hzRuAlSdqMsDz7SfoVKQfWUGN07SpJJk5m
0XXQvHiZISNGdyHO+OGeVRJyLgkv/FK517qNqjtrmac//azT8am41CV45weP4zVynyfd9M1ir8mm
gci6TjQS6THJKC6v3HIMm8mQIOdxsYRhgzJdIBq26gKMgGlt4XWpZbxcq3soD+1/tMmgqOhkSgjN
wx5YszeCRHjK5DvyfcGKrCFxMPhJCcvisKUXDhIuXBpcRGLz9AaCMkVFmj9q4f6NDlrE4s61MccQ
FBrDlrFmC3RlasHNxIMZHz7Mdz5J7D7YuU6Bb5oqb4dI+X38fQNU3+IK06akTjTFscsKfqI6hqu3
XcZFtLzLBz70eVoNKNQhcYDHq/hnnhhaad+mWZCyy7/yBCKmzfj04a67H7DW0L3c2ASUGeP9uLp2
uKUbJbz4HE6cw2mg8Wu7QYEGMn9b2nAwp+g5chJ+mKd5gVUSA4bVMsdsGD5T3MSXiR2tBi2MzIXW
xzqn08j8k4rhcf26Wc583oGZx44jrtIymIG2vaZo3oL4AmlN814YDHhv0DyLQvNPOUJTkITxWhth
wzBocu8G5Z4+aCJrnDjTdKyG26+hb8eI6Y/ITHdqP/rO/6fGxhuAEPetq7/rsT9HJ57ucLS8RbH7
0ebbcPNtdagxv1qldgxVbOUONR2n0o38M4njM3GQIQO7WHo1D6OzTpdfsrIOxk/1dvwR6/Em9WCZ
/9OpV1bEA5IulgNpWF1jXixkco7crfPHJlJfENTpnLu+reOM4Ui/So8R02wPGv1qvOuL5M8d+UPn
pnRZSgkiXMhgQcWw3oCffIMpvTcjYMAtTTb4yCmupgeLIsUV9Ndy+YM/Oc5UYc1TXD3lzb7xmLWa
idw9QBuykG+PPBHj5rZZiYNv5NdFfzkCb3gZZ5h2MdjqkgM/bgkdeJVkapXgToT/C2PuTT2YO8MR
mx+Xlw6SvHWQqi5Sd1jcrU0vOOd6kZuF8qMhLAPTp5ts8V/OUPdGlARaTotZcI03lJc73NVQfLGl
Awe+F6yNxh+5Ly6LZql1RD5OahHKDTu/3QEatmE0KO8fMlJHQvqzWXKg/V+blU21jkbsLFoQHo1g
Pmg3p+Dt06KofXHjDm53KoEMLQC4jgE4h9qyaYw7chaaeRz45a+ta+P0ZAAln5ilggum2QG5Sm4G
woP0+UHHw3v3CfD1s2vAk1hM1VfQ++ev2e1Q9JW206y6/t5ErHHckAxHMykVANUBp3rZo/UEmlSW
MIAwF6xdSURgPLzrJQpGTo6kKnTYQm5YL8djjkO5zKMH1EbAtoflwy0d9aX23zFW6g48iAQWePuz
G05WcOb9Ktq0QT0E+h5Dscqkq+gWft7jmQ3S/obqOiKGucAPq2MgRIpUvct69Trlt6oV334uim9U
yVHIU1WlajU4ZiT671XapoHx2bm2I8pLOA7cNiEUMk1/dn5PfhF1BFi85+SkfpNDrEr3rq+mtho9
cnYwNLBO5bw5ZPOxGf+9YJcxqmCu1LZw8mN+C2ENuLQoI8PmnftYzrTQXw2Drpdp5GlxR7HsWT9K
CZJbQWR8Awa0zrbd9Wv6w4XIP7NRLlZZ7M44z+Cg9KjsLL6ZCWI2GxnCAU0Dek+GoXq9lgXZooDD
FqVVfJcdXZT/Nk3TaWYJP1oCOmdst15nubcYEnWjZxi19iAhy7N7sjDE3WGdrr9vcTtDBCHwVjGp
dk3vYWmCSufoVYS2Ufz4V0+I9zbkEBv4KR3xQ/JSU3n1fsAKqXh9GDqb8qZkvspISknby/NdkSzZ
2BCvpGaDXvQwzp0curogS/ntbgAnW+ssUdkYnAlpvpGDncsK6uyBVqe4TQcrUpfihbi0CIGknUSH
mcqwL5BuxXv78/A+y3kYirLuFDT0t4if7yKZ07To51K1EQQMM/n7KYmqyX+jzYJOjXLnDLHP2BYU
XYxbwnvHGkFF4AhZt3zMRKQnRZjRfrkwrTayqugM5f/Rd3oVxIXyDKqJEY6Zjk/J66SzXGCE0UhG
V/gw05FM1lW38mJePQzJiLb00Rz4mdcSGRuuE3KdBjlT2UuD+qHbo5ukz+nOAUb/ekI7gSj2zMKd
BgXYOX5Kfn3+XDyi+yQ5s+b+LS1ul/4xvWQM/aoryKC3LbF784PVeleX2uzLw/s99RxAGiIE3CrK
i9pkXma0nYEXrJ+AriDN2K3RmaoyLbedjY1A8SWNAzgFJqPVuIs+1IeyHRgMog0jBa2A3hotiNXW
4mWJRQPK3KpEvcUeOrDtQsc0wex03NF8/JEE8lTh/r4p7377b+yagAiUWWFxQrVHJYNtcXVZdNaN
WzsQFOc3pKV9QfUD7Mx7gKsMUaLY4dnngIqXBWA8E4ONKuXMJdOX9k68+3WP2iYgyBV1Yb1S0mWi
ktxHI/kVmqKjubg8V21qgTiTPYaP7JlSvLLOJsd6nSnRpOgAjL6ivNjgosRqtKJyTapzfZM+L43h
YGy0h2fqq3/UEVoSWQaa1eFasGDERu/UY+/9LvKBDsDMR2gPTnGjKYC3oU9GUJzfucfdmt/wN/YU
CnG76TGMcGIEq947k7KrB/r4bzzAg/zAa968BQsIoqlAxE1UuGcLgjSm0tdw7NZusqV7Ai0vqZrK
nyOvYdClohxu0k9iQjrvn8uvABGBNs8vF97fB/mrdOH+Egcso/7ItEpjg7L7lG2QEtmB4Zt/ui5E
s/jNxB9cYee9RAeVGgkI9f7ZH1oxHechvUqoDqLeOOWHB1N+3ODSpgRhU5a/k9d3PVVDJoUJrD/g
yXzgYo1UFFId5fZDjf1+uUMawdG/f9fI9FPWaNOh1ZTDaBpYcVokQKUEKpuKp18y+46Tmb8WkRaa
y6lY9dOG9uaUVoNCa3Dvkj/ZKcBoiLcjfSmAnNdkNnHAlurxxGeFGoPhzDOtCbjIs/KTU4A87STF
UNHXuZtwxXoieVjpL79+Tx1VeAMubzJT5CXxlG4Y8dnZRQgI2KKejt/Y8bJ5fOu5nhh/BjdBvYxG
iAtxExHsq1qiVLpmMIEPMxaxJOri8VLFQKAiKbMJQg/xc9vT+RtxFIT2J2gDNKaDzrl03HEQ0JuD
agHX5SWJ6YMNbtNx1XLrmipR75QPKAC3IlMgVpcAFdc00ftyPi/v5wZGEgnbRq6XdmUBVPutYlzy
BBc/iSyZ3Da4OjLpUuZXRkXLDTpGjYnPDVmLPKzraB8QP0W+qKF0Cgc1AOY15gOqhhnTD2Fi4mIs
VFtz+KKNxUPMizkt1ofSf40bV7+fUX4CBgwKajBZhl+xE/OSdTl5DZcwStUju57gwx9qnJ8hBANZ
0zwZ0jeI3tq0lxuR4B2xXThKcjMDVH/ieT1DvD4fJWmVwz/it1nEQi03xGQ9WFevdkTXtiqOFWbS
1wcUNXiqkLEFjk3JAgZf07VcD/cx/K8f+3W8MvnKUsK/3zaOOGq0IWDgiJWcz1xXvrYwoRpI2qJ/
/6o+l/O1E9hjjbnAZcX2Gvn+1OTBPDsMscPyOOyMfFndP3pWh2eDbvULH/g5rvZ0mAHI9Ec9t5mu
5gaKLPQA8+xdo4NfJFfyjKqc6HL570B6sedV+KpFA9peIxPQZwS+c/UQTCHzV/w+qmz1PqhvIo/V
D6GaDEaUj7mSZJGFbdF9x1vz8dx9VwJ2/Rknw4Kz5CRZsnZn0fEc93TwKVKe+2A31UGW8Lx3ulK7
P/gb+uz6Jjrxggs79HgrsAdN47iTAlKGY8LS+fjYRCDlB85qEN6/NHPx0x5D31EYW0OmSC7vJQTK
IO/XhXv2vRAWBzAWJy9mc745Pp5tM/F+oIPM3D3y0AcxkYd4MDOh28+QjkmsO0peock2BNn7i5Fw
hfx3NYU4oRtEMNNe03biE47aADqUDMqWLg4QfBABJkVvw8d2TuT+Na5Qyov/RF/uOK4whyf0hXU1
LaQFKaSCxWsHQ1RD4sijjnf7L6Q8EpKSFt3PrmZurgIfaqKYCHXCSIpP4007XdLpfU+TtweAaH2G
bjaxlwDBDp9qRkTtdcYinlOthWoRfCfcVOxt9JrbekQIg3BnA2cvAF50ElX6LgXvoLWntVhTdMit
rqgzfJ5mN6f3wcAk8VxruWuvCLKmaAkhutDhrQ/GgERsxBLg/GFcr3pLtbLOsHzKATi1cCnXyLho
RV1qvdfgkIh76SbVSKzMk+HjEnQ0PuWpowgkziMwCZMg4bLnNfdmpzQOHebyeutdECJ+u3IXyZSN
fQcy5KFMxcZuEfA1cmv/8xXuem7G6Yl5uwFHsBYDD+psYUWYv7+caV1eXd9d5f86b+xfTXvpqZfP
5VDHF0oWU/adJHuRtLyBw1zzhoup0jRv7UaWGte270VxAt4Mm4bGXHf1xoXTZMxJJ39iGIs4IsIo
6WYLA5QA5qWiD7sFcoNAecVgg/ajwdG9XsDJCZZVQsIJVeI8BRC32afyJrvJRuJe5DJs/8p6IAwC
iWPuQemDtUZO+joDDxvXaM9fN0ecgJJl2ZcXeARWzLdEA9vNoGrdpAIFsi6P+xrlvrIbNsJaJe+/
YMb16x5ARcXIHj6D7aNHaIiUcqEDNbyf+ZBjEK6ylAHVqHvSHe61a7yTu6Q5gmaiNXJz7zPi33cR
0i9GgT6MHvIa0Lj9JxGjAE3SlIBxtfoOJfHZfZI5uowW1RDybr53orJSdFy4edGz/wnZBVXwQ2fD
aupUOHSTk9MEFvV14LWQcGn0xMhWzjZqy2J2TuETAjbc52lWdeHt7DnREdoUtqyXg3JhMhYjNQE0
TohT80fVtOBRgdhbU/BuOUChB5U1SxajUJpbvJOM14zpMqqJoU/8MXCL0TY1fGk8pP4y/Pi2UA/J
UkAjo+SdpxmGcxeBatoTwE11jy0NKMgfZyPXygPPMGKSKr0XFqcsei5sGqysbtLpHTXoIZx9kpPn
z515qVcDs8KzIYAcODss4ny94qwgNvU8F1XqszDRL/HUvZb4GPYFeAkNKMXUqJQRbMxtXWkiRz6w
aJzu7VgBVS97yXhonDOhAd2ZDl98kIp7zCYJbCUKNIiErtjGwYbn5CPIZY1wVb4ZQvLgAMsOPg55
xSjfCA+scNgaFp0fAUuJQlKh6oydpWsk4euBoLT1X/nH9WErLupwR0kk1viQKJC///fEs7VVMkEf
Ql5+WFwpyTa9RoGD3A1yLez/CVY5T+/nTb+uuuncWxVMjjxAk6pdm6pKsj/eLKnljQU4nd1NYZuz
DpvVqADtb9GPKulwj8TTzXdpi/JIGjhFZDnV6MsKBNXkLGNM87ewPqv+qaGvT+1CAw0mcobb+1gi
huyltHEmotNZ9T5xGGm0grX1rHM1yOL5Z+eyVksIhQhcDdDip30QwEMqzJeobrUbIm5QcaRTCvX3
K7B8nUAL3oao5Ay/cysLsbM64/V3eYbzB6JfSUMoMFq+IXZSXHGTQ3Zv2XHVnNajC0CerlzTsQCv
ke9kj/fOdfgJ0/zb6wKNdyvh6DlUYgMGWOyJ18UQHmM/oh9S+pAtsXPcVd+RhJUv82TAMMq230w3
UYpVjD5AGoQsNxv5I8lUfr69vVZJ5y84WjrBV1LgK1Cb1zDY0tRKwCcB+X5H22zw2ITsScRTJ2v1
F04RJXWM3pMUCAoP1M0bq0lH9ZiMtZ4R3YuTNPGgUvjWrcdUdpQg+2ry506xKnUS2qNWGfWpAgIt
AbvAG+OZwWQcfbhhZLpLSQa54iOrbd6KvXy+xrZWeX5hXILRpTAF0TnyiC6KxcpMEItREVbnFIVg
rK+KbBxtsYPwk9iGNN5YNrIfBXG1IpNtvrD8TQEDnqEKP21Avi4qE1STSafHKycMyYGJG6jGGjM0
AVHvocSFVnoTOutKnLFLmv5h6YzPvaLPnuYviM1ir2kg/4rfpVYQvYjqoXxYbOQlvBNuXwBxyGD+
WeV5/Xd0eop9Bwg/nODx9IeuDRcMSEV3mEMDGjOSN3owSM9hFPXRqvxI5/+OvUrpiM8ygXRd6Ovu
ryLmdI9u0aJbMNDQOAzp/NymkzB58AHW3sb0d8X6EwykDAPzZienv4qwgPJhFCkJgQeLa/ZUnrFi
mJQxKo1rkqwvsMKpvBDXbq33kdYqXM5DmufCN6a9spFNgFaPHNMWGkcjuGmRtJrOKCvEvWE2m5vr
avIiKddfEmKtoedDNryVV+Vigpu4XFagO1K8bUYJ8RtRtai5o1VkiA5SEDf+QPo29V0LFWdHznQE
n1hRUcyBMdmiLh5JDWb3qEehEGPBzImSNcSdkk4gZI/lJvXIoSmPuP2M5CuXWsBv+DdnihJFbVZH
5VIZNuxdsQoRv2yVLFe+kzD4C7DfX4yPc59QkAlMEpP6Gw40U9Cb66/05tInAPuc6dHqKA+riniW
9tC6ZN2nuAkYfYOlmDycwss8cDnNw+MY5PZhbbyv3A4KSKGFIQzVc+dC9F9LOrYD28dMGa468Twd
XsIPNDqnOPgIOg3pV1fveZ8FJlcTCF1x4VDKu5f62fmMuQel6rxgwSfhyahYVPGkm1Z9/3yZiWjh
urzhMJBH2X0DrOMJZi5TneHV+c99qU0H1L1WQzQGEJLN6ZtNk3yZWKPpph8bZXnsExu+52NQ27yK
8Zoe3v3nSSQ9ZfrqXxOm/1iIbkSJlDMWMpzTAo6tr/ZndsAT4lHdNf4VqMRBz90kB0kyTxnz62RY
Oyx/Kx6IzIStSxSz2G8JQGhhk/CRbOeRuxCtaOdPFF6Ve9xvRdyYquao2Q4Cr+2KOyuelNP0NdS/
TQ1P2kxGlVfyoDjt3i0/MyB8zXH3wF1cHf7b4c5rnTh+T0bYTUWwaL2PjCFvQ1OWgUweRO12KHiU
fnRkXocONBo0t8Mq75wyY0GOVxyuMDfigMzlRbhbwT3rR4x0oMRTqkCIuguY4ZJkS3kfYJVvFbrG
p4ck9r/4qBgq92BnmCARz0kbjl2zO3GgBid0Sq7oXXofJCwz/9vgmhIww5orJes+TQesAOqN1QzD
k/QkGAc6mrmFkTDs69AFR4gONRoxX9mGJAodwzKRGnRfEj3OLeArtuGYHbXyO1RgUtZNAWPjfflj
B3PXwc8ZK4IM9g/1QCW9XvXHKrIAV2GN+jnpmTTUMuuUgN6GyKGx4jTTVOtqTYmNg39KXyrlIfUV
qqwGiRExFk55/BCh2xHQCwrRHmtXey9Dn5BcDdW7flng7ioKF+V9u3+wrb5f6H0VHLIEnC4RRBWB
W9zLoYByldLj+/ye002JF/rp8lkGrO/cJPe7b+q+tH8C6dp1N78Mdem+RyF0odQAXANdmsSqd1Ow
USBVrIuzO/C1SraZ/AmcmgtSyyNOSMrT2vCkstVox0ojrXAqX5K6DtFLPzjieOdiCnQAZ1dLHzH+
+hA8gJ5LG7OTjeTJcNGO4qp7MP+xgYjgT0mBPuDiQSdjfBCeo5FMyLmz/OEi3W6hmcEdQaKWPafE
BL7XaEhahzRNruuKvfQkNuWWlJDDeRsbXzkl+kDzNsu3/GyWRObywuNqi+M+0jatUpaelXWvGG8F
QxSkkad1CcigkxN0QX0SRA326+RHNWigUNDg9R3gtuR4yTWtRTb7QlJr3qlui36wJjUwBzAxR/Gz
w/e7hfctjUonm9wul5VKYCvhz42B1Ze+x9dvba/VHlMb4huGXK3SJ04JvkSt1oIGhUP5jNq1rhmS
r96+kTnWK8KXeCLcrdyKJe5o5aoNurbRQ4qeeJvR9JVsdfMx/x7MLjT+szNMbL5exhpJwfwiSSmH
4c5vSiFo/L+hL9l34MxXeF6Ad/7tLLHQnxDZ1BoTvktPfPA1UkKcAqoIOYByKyooUA28nHEAfuIc
YaK0Md7HYvghSSvDbNGYBNTP7JKfMLzbsisvyJuFKPHyCReAC1H9lT7W0fFPh2QOBDSTGkBuq4Gu
Ov3h7ZN6PRC8XLGZRkLzWF1RGJKvpONNXyYCLPGM3aoo6VHtGtrixTw9yaYJTUQgMMpcX3MsbJwO
nFuNQjbxtuo3tpXQxqNywzs93WmnwjyWxAO6UmH5SeuhKB2Zkfoigf9MsbVnwnJ1PhEPvkhaDnNC
ufwnQxzhGxCaZjZQ5YGlp4J7H3Uo5EXi6RDWk+q5GMz5E6klwbn201xHM6hdwVKjg0hDc2Adc7eD
gEbRHtc2jEWdp462LaS5d5USe7Qtf4LNvKGPCAeBNl2YblCPbg7pYmQ602iF9H1C2EddWDNEprmD
jxq+rYseHa8wmG5lWRymwCtIX5uqobfIIE/YZqBYIOICAWrlhzkdMMacojRM/dz3ljA+gSitmQ9x
obF3EfIDE86oMfERLDjkUUjDLMy1Wwwn5lOCgOWFs8IouEoPU4LzV6l665ahn0INRHcOz4w6WBxA
FY59mEdh+IbwQtDt3h4NyJ7QR6LjI+M2QPK9wUUKqLO6yT8YhUmyjBGXxOfSIbQR3wLItxwnui/S
wE0a0skRkMH3BwzgVPJtXRDI/b5XDwEpqA7ERYupyk4qZObErfksHK9xFXXao3kpTVR6/zrgxrsf
UV67uIhU7KttLA/av6RmiDSuJPAG4sItHDIbMLSqUma1NC7jQY0MBr+xOuYFHIIMkdvRVo5Ui3d0
3Tx28LLN4jnGY/fdjBkkuxi/WJkzbnPGO7HG9O8u+xsamnOtCzl3aPA3jsvYkKstnjU1EXa+3jV6
7IHK8DdtIuJjkNokpku1qsfJNgv+3xVVN5VVf7jWQFIrqLzKCLsLLII6cs7Yaf0xvdbLW+7HY+Q4
lOVo6QrSIuZJrLzIIveAk+p/mSS0IZ4k1/5vhKuV+vqufs9ZwxM3sGm+Jx3EuxoU+lTr/8LdZNP6
Hwn/OPBOsSLKHNOOdxxGi8uS6uAGlPWXRCbZzdSBK1GC2S2ht4yS1aYAHVYY9Pzv1lyOWas7IRmI
FL5T5c8u4mE2DcMPjeADq9hqF4hV0wNy/2diGeOUjuhzwKM4O6VqKcMMab1DYDWr+crZ/7oVK5GV
C1mXJTVsprT9Z51deWxim+GPw8ritOM76arzMLwghdPvM1yaMmLkSKV7jNSAQGJv1H4BUkvrzZwV
UfH6GOggnXMftcMa4M/3MzA5LiRzJnzDH9qm96Fdqjb4t0A7nHleshOajH+GL9ZoW1lRUmCSfYib
4UXPttHtoZ4c+SJXLuKgivvqDVP7A8C8iuCQ9PrIrunfc0zrlF8VN96jPmHV2S287h3PkE8kFoQU
ScyEWh1Eu9mkm0kTDT1Tr/Nzg6SaRzOG2WS75qTN/hwCvXYo+R6WYWwt7U1Nsjf/2hLUPasybWDD
fhQ5fkuuX7G20m5QzkTcgR5kA2DFs1IeQ1apOzQJIQ1e4E1FVdll1QbdsfZI5oy/riXO/nLQLmIk
ZqhfQe1CJE/xDQT2WNL+dmhoTq26jhSkB78SVYlK3JQHmZ5pSxfYki8pXRrUbRreTEHKcGkLACpe
crlurkR0qmgGxYEzxZtYTGo7uumMrFwt6pZkXiDprkjA8tPJPKpiLunpSYjIZlB1NXd2Fvc5X1hn
G4aT7rr+HnH6Jbck18Zqs/Ywmj5U3bzeB8TK/swDPQCp1mxk5IpiGoNzyEZVONTcmM2NJ5aB8n5x
6+oT4ahary8oIqU0ODeDUDIcSQVRHiSj+Gd3d2twig4LSPobOIqX7gx25RUNBkHn+UEOzJDVwiFp
InDUXKfbKXv7Qfqc0pUfKZl9VsDiIyIR2pyfXyV+D7pE3cGexsCzgw3nNoyd0RRTY0kVkQJnd3Ld
KPdg/AJddSPFZBbmVtPWBJH260wYAoUbcWldSx/jgQKfL/6vS40uB7RJamddC8VmMc7Vg7atDsd2
2Hb9zFxpZoCTfLpru+CP6j20GBQFbBUK1CkRgNbDDNBSsGsP6YfiR0Yh60n7InwojTe5W5epK5Hd
OZwy0n7EGp+tOgpx405oI0nfdJNry//RYfWgHAfZf/kMQw/kolOlOXX3wuI4PcwCxEDh9XuyYjKy
TqFApESmk6h4vZZny4kVUfXxaakObir9EzcCRchgYdXiSjNr+fTCauuZrZhQOBp+4wE7tz9QjhJg
LIlLrZ2wvoWxx27jVXo7EpWk4Y8L7Vb3vtpUOg8i++21BjUjRXkTVC9h4MA0O/8wfv4V3wamOR8d
1OZZaOvF7FSxPAk69suioo6pARynYjESicE2Fiy91U1XjJVBIgxH1k0hxfiitI8580IowkW5JxHQ
SAqGLhRHSZIHPoXcF1dSo5909riieU+iFHRI5GD5Bu0CyIBm5TRlM/SLIoYeshwa9uuLhp6BCyii
Q9MC2E1itHkkNpgK51LlqjCdghihAw22msMQWAx0ZYMjv8m53TcOcaDhkDcDe9QEQqOFPF10km83
MDL9QXEnjhd3tLdSNh5MEDWYcXTwKFqrjL4nPkRac2YwMwLRAAeC2VSxv/oB9fWM9o4+sYTnhl7C
srKfI4ofmqGAZzRPwXdMbYaIUUftac1qvb8oRLHhsVb3HC/ea2tF7LKE4biVmb7nUgu9MvzNgdBI
fUbMDOOZqgpH20CufUZQCLDPEVdDnWI10sB2xxcPgvHsO98jKDa/GJ5m5/PZwd9UsVdxGUNSFRY1
TPCEkZBW5u/ABERAYlLzUwjC/59Nr8HanvsTLH79PwPf6k0AdTF3tAzPKmqqhDlpxw3ydEvNlZVk
qc32GcspKaexQJlXVxk1SLB1weQXn6tiIscgXvwXvT8JIj9pNM2Q9n5KY/iRhYnTc7iRGaEROEEO
62QgGV0OC/+WP5oDsNXhKQ0pRBbFITXXSVzvjBKZob/KCXty+cwujct15IkWQUDmtZ2yUGW84/E1
zP9cdwZOUnsLSDUU5SHIZbghIjCzX2sSG5ziVmg9Zr5+sTwj0wPRTWQbuSb6+/MgiZA4iTauZStr
BAP5IEUsqRX3rZWwdwMOgovV4azQs3i524Y1g+a3IBWO+HxJDEYmL4Nr/LNvTmUl9Tuyb4x2u9qu
b1B8FxKtlbQ2YjTzZcbe5AX4WA7/832EKJwe1uCzOWiqaHpVc4o+BjVkJtaC5TsTeJuhBOANEVtF
qq17kbn3pxSzFs8WfRTWnh62rBn2Q7BPYMpgtVRxxxNRVNW0zZsguSDiHJy7C73oyw+8jk8py9lg
Qhrx+I58qvGIGUUVFbYUcHp42vzcS7kqAqInALsN/wfBlykxkKTgn5cDokZIX9VtEsd7c2irz0l0
V6h8ZoGX1T4NOnsdmTSZV0PuXxMSjy523i4/11Smy661E63TF+osiUScPNdmmrFiDNQPWgili6A0
D+loOfa1tdA+GLde2KTgXSRfYZd7r0kiiooHf8L+++70EExzrGfR3V8F7JAeFv84U+TZQ0FX7gWS
o0E3+0RFgFoc18GkIF/tpNCJ1gL+AYB/41S4mRx0Y9DTinJ8l4ZbSkPIOg0W5v8rOwDTT0vbGwHr
1N5i3NPaJLsSzDCp5GK9QeUvsyqFTCHJ1W4uPin4dT9b9ZuHhSeDWAoVlbI7wIaeRAqr85w+SL6U
NC0Scmq7FyWVq9GmebCuTIp65kEiA0KZo5JL2NJCZDd7og9ugZc+k3hnCRe1I5z1rqTnkRTD0NGQ
UkfTDGjpZgrs6TIMRuuuOiog8qWgnVO+YNKZyJIdZaDj+8MWVr6WSDIZKqd0JzXsg+A5RsA2uMs/
ofhQ5VoU6O65piwL9419RNOK/65zkTgLhN4X6v32zIs8Xwh9Be9/YgMeDjBKyEdxgo2ZHBqiKoXv
vqI6t7lrIhEyTWIkf6Ykp1fHpwX793YYV2tHLeT0vKvsfCWR+P7fvkgTt8qWDf6R/oEwFGQKo8xy
MlxNYsTw7UmojKD5KN0jZmDZYSHfb8FNkZqO4ab4hthqdxjWz3puLaH0UFa1G2j3WvspH15Ir0nx
PqRAYUJ270uBGfZowrOlOdCdibk7Wy2z6dFYiEMGVPCdW9szNyKgdBgTowI2EdbSJzvauUQBPbLV
1RbYsvrvWuqJv5v+Y95Ch3J0Z0VW4e56ewogjPjUFH9V3o8ofdEma/iJutC37uBEBugGLPyMXtaM
KoOlUMvq0ga2cJH5c+QUR5SqvksjaYe0nneXzxukgyUxpCW+tg5O5DdtbceHmud/ckbsQEimaFhj
gxpBUK4/tPsBTpgSpI1hggz6dKj/xNgT7w/4/Y062LbcSqCya4k/xLiEborWdada5QezVhD5jS4S
yvjmrK/aGlKU9sBAch+9iQf4nnteOE3UK3CQNEVUi5hMWoVtmR0Tb98CQSoAlgfzuKWdQEkN5Y08
KGSG7RCIl1Zwa/fpnXs/RTNiBxosld+yPXKJc7g8Pj5jkFtKgyqLRfMTGhd9Rz1cddtan9pQVxw0
x08DWD07uHckUi4WQuCXITuogotVttBGlSF/QdOlzZf9P0Oom3RUZtHKBR+M8hskVcAx1c86b+GE
XVguiykkc85Qapzi9FsQlI0Q5OtTw+/70xgDFt5Ubfs+H0ia356q4AvpqWyoY9vNPjp2Zp5Z3sdp
GYcja+1r9t07/GgC3HPfnxca1YzWd+7/67OeVpvE6Hz56WpBiJMVHDcyMeMKLfrMYa5ckRAUvFn0
pbi0nC1e6P7i3WqaRwunVEb7CVA4E9k3JCF5J9Z1vOOgoZZY6bhNXqjJVQKJA/r6ynfbCiQT70NF
/QalH6ZgufF1axZNhicpQjhIvyxyTuYauI0iqTTzea5Ze0/H0Ti2VbQpu5UP7IfNuvh7u23fAW1e
b6Me2S3s39yRLlhiHzzhlqlgziYzTJUzk4owYl5bglmHaYhTtd0iUOgFdsLonjALZJP+O5BLovpO
7V/0TTKYwPF5gCTjfe2kDpyLY8aijaYkCMWuAhLCvluJc5ROYHsTMiQv8nRC7IrvUt9BV53Uhtvg
nNnF0M7iUGd5wdGvd7XcVNQqT+ZsvUbyo5vk1rVsfEyOGyv+NbuHVA7OAtBb+hsdBhFLa2299h6y
dmXtnCEN2Bm3A6NOokWBGOnVz7DcqgIMrWtgtKv/jGA4rpKadczC3kYogPtDnu0yw3ig03iba7G5
LPz3pxhdaDezEmzr6GViViBNYNYluNB+MCQ5MmYfKiCF9uabnVzJy4ou8XAbEq2NHLT2GF78OSqZ
9AHle42A2nxclIhsFPYnmQ35dEot82LlvCIHCkdtqkQ6mKZkbYAtMrZLoChDvzM5+zNMDg2Byx6X
V7okNlc/OWE9MGkGb3QdoAuZVt/Eq77tVQwDEybW4Yftx3znev7XBz5UTeaHgegQKjXSzIlaBTxN
uvyUx7e+RrS834q8myKt21PAlQ7BRjE6wbMmDl0D3uBvLmZXmFZHD8WEZ6hBuq/lqodlO0hMvr4y
LHZjt86sYwrpShqHpvBv3IrKiayqimVLLLY/zTFAjZVzy8sNvRwWXIrwa4SExkFheqZ1JIBhHQoX
KjrWBA+kW/dmH24vRJstgvJpuDI0f19nFZOuu7dsSdOSCcGLt1A8GR29wQoEDIt4b8ZJRS3gW/Ei
SO6xK3oN+rBku2k8p8a+aSWKJHUo75wXSHLPVAhHSS0CG7sZzGxN18iBnPJYlLng7IQNVI3Ppk6j
oDlpF4P4Vf8IlguyIaHLVs+LrAWDaEfxaV+opj2pf77D0FyRhWLKd55QoQasW8Ul8xp5lxkzDZxf
j7Isls0JRhQ2265GLitY8M7e3j/8m//CSfIY1lythaF/+egeEoq1rYWdsIp6WVYeL63nDQIO0apb
f3LlEbzKVP5N247PAKwr+CXVkZLp2ayEMZsN4gr+0BwgrIcq6ucHmaQ2iKWUHmfelmSKC35A4pis
7NEmp+Jc1fqcR9+v4WUFXF+pHZ3vOtkY9frM4HRb0QI+J4ymTCfXuKtv82a+9kPrYSCPFBVRO7Ya
0z45pp7+e1+y8A5SDMUM6vBF3BBdbTjJ40/0vA8y+Fs9TpGqpyuX145hHSf212qa9kWgH5udzXcg
WSZqiRnk2s7WLOFowOWhoyh1ffqALkF2EyGRchHR3ToQiUnjCHuEkIc0qwSOcMeNkpbklnK/X2b6
AG9j97k6AM8ofP83Y/3l28V3R3mi3Va2/gM3oMj5eDWLnNpdWFgfNDPvQIBknFiIb8ir8CvJ06oZ
ZqXGEbLQERHaZoRbO3MfQ0LGeW+o25M3qenzJH/ZrB6QeoUhFKp58W6KrFXApSYpebxgzUdN7l3p
RmY9UwHpoMWlDyFHDHnak3CsrmdyWMd0sD3infNkceNu8bwY9hSCKrrkHgpq7NRwE5FN8+ZsLvOg
GvumuG8YY/0l/hfE0zpMKjyIIyJ8fWpkPrp8aqdNSWwF5cLPbTj0t8ikcKegI3qwVV3NLFUq/02N
00AO3eQjcZ0DVSPeTU9seSzbNdVuV2X9GuFg0UBgAiX30eWD6X9lHcwFPg27zRP1oqtIjPIISXtG
yB7rrXJsNLyPVfE0si4LxpcwPANbTwOaK4zO0Dn6om2bAz2s6VNPXVxepFWqtH2+8Tanbn2QcwjG
Vgl8LhsBpDAw00TViTs+whd78nZX0b1+HFmqvlvUk6d3uR5EUvsWaCOXgoXKt8rQvRKDvN3vSUsP
felN/2aQA/ChawblMaubYG2R/SksTegTrHEP3SgSHNWsZohY/68bDwaV4E9tCMWzb9wooKYK8kSg
M4SiaxaWnn+bpuMHFVcNNHHJ2f7z/EvpWDUoVk8GXZfdqSF3KWuOBYOy97D2F0Rovr8vUYhS/cV+
9YsUDGTKVzk1KlRZKcIme3DbbYBV9u3r03Qo1supwSOoPDFXby6JPtVxkBKjMJhpEHIBFZAb2i0s
y+rnN6qNaMQ8fxK43RSIWfCCttVnyiXgLUhGnuo/mNocy+cMH1ncuA6eNluL6m7p/oQ3bc6t4V5r
PuS+ZrqYp3lxaZMUWdDHidlMrfkAK8udc2X/JvHttOssMpEnM16HYc9YqyZf+3dRl65h3GuB998Z
GHT3TA97fjrhnri2sMtxtkUPDd/pvmg+uihxUJ+hN3ZndHR5Esc/uRHAY04RehFJ6BIR+h5Oo34M
9Uq7ocUBbGYPPT80T3JNektJAcBrwalvQpP5IlctiZdzSXDWsxJ/Drk0elMxZVEPiEheaUbMQixv
8n7h19osX1D6b8aQbJc6H+z6j53YqFQHuylNi6Wkv6+mNbVMHdqopbcXLEP5rFtu/dxPpbg9Toaw
iFlClWk4UijiQRWadvLdnBZVRYPEORyIRo44vC6y01UXVQNeAdcoyqWQBC/qon/rJYdb4kxIdyM+
N4Qs0OpxzYmh67kQt2uY0wYwPhUgJ3KSrUkdr7ppY16iggWytyrCpt2scRAVSCHDkNgCXdogMqb1
iYNjZ8KpvZxxv9z53uobCR1YPlPixaAebpAzQXeQ6fzggO3BGR1+B+lLQHaPYaXaYdav0OYp5MM4
9bqXmTjnbKb8s67gi8cFhNQkk8itzeJ4xDXE+mQQl733ElRmnEJ7DDLhGkF439iqEsmISThULPaW
If/WgTbrrADevoI3LlV7SxfyG8KbKuX4Gz6TQWf7zOzAOPqcSrrRV90KAwsgb+EV1Fvo0vzx51Lg
rQspdurwtROMPF1CecJe93We24CE/jTxi2gfDORo7H/05mWYs1wI7F8BviFDcDz2lVFvv7XrfL23
jimFMh46awnjGz5rsoLfwYEG2jWIwyEJ+iLkXy0/Tlw2FaS8uG9uiuWpibQ5bARi6YKj1ZSVKUvL
w50XMjNULPSbxVkHTZnUolluDIQHQUFiCkSBV0hzLN4Cng4i04/2KrTlqQSjww8eBvXujCwDmNp5
HvelDBakjewxfhFIoi1NvZaCJJCFiqiM8z1AGMVOsnQynP2VD6BNYsRuVIJeEGyhQV146MqPDo38
/nACgxFwmhlkREl3yfUORmzvPk0fH7mZQeKvFywiG2tWItGATEy2ceD+rwfLHb+4c8xcb80P8olY
5mXSQ8XGBDvSHKf4n84k+kkBB2LgyqPB9ToWSpt/VBxhKMeQzRB9yxJ/EsdOSu/LnoDbuMCPENQi
YTGi7T6we1Dr6L5wGcpiTyiQjlSbLZF6PqmgtZGcpOCKOAqHZB4rY+zge5EtFLcIsBCpv12JI0bx
FGrFuFlLN/2mbMZNk9i6fSJpzN+L3FKuB3hu94XskSyd6QWfhPZGOSIE6NehRKHylrbGKBO3Y6KO
K4/f9TQSzFjCemoV703V/xp7xTSI+iw/1+/nacqITlCZgwfmaien64mJVn4XtLsTDY5bIGuHMjuW
pgRUUyboFoRM4TKnr8+GJNZX+nv2EkxVP4gp7ny/ioDoMcMECajw65jqafUVD1PWhKWJGs9tkSzk
sHwd9POXu8JPqdnJRhEL5s91i1IZCD/tix2W60DZAkyUz5cNACUXsusKkxgcxtUnr5Q9SXj4zGoS
x2FCuv/aWfbW3v0DPzWtwE6GMh/S4JogFSP28dN4H6VPcgJuHMxtjbd/PlN5nMxt6xWtw1+jcKvG
hiYcx0SXNVIwxj4BqVaflBkWl+C1d191z9Qqcetv1gnHmkXbpdMlfPeIgsKVkTnuPLGf6Lf+s0lZ
9OObg6Pbir0p+1Dw5dmNNy0frPXEYFYSKNcZi7u2kZDIHDB1ie3Uz1rEkAhudG1J2wq6MDVan/uK
Ji0v/96A9v7vTQL5xiMaLNXTMymVcv/A9K5GNlMdWeCIqBMedbKdlYelhLy3W20d/ZmNHhEvnPdb
BAHiCDnkWZxIP4MYIRSGTKKTTeRibaSKK6mQMv9Wpqg5LODgJb9AZ6T7z8n6FKTFsuoG10+6R5JI
YnIBA1mSCPr9F6dZzQvjMHiBq9Pd6EYbnb+ZGx/uXw1uwWzKD7UhvTS2QdXW9MdGWWQ5eoGdRbmM
2ttPQlr82q97huiPn2pmasmvIr0u4MQn3uLluM4SobN7pV31joVrITrwCG6GM02B4GguwUmtyNcH
y+yR0HEQWru5jNlFlS5H5TI0lW++iZ9uWMaAInZ5/Xfby0R9MDxYV/Wi67Vy+l+HW6glcnIkfeFC
nKhyAWKpglgf1+nl8hChsvQ1cdrrAjVE4mF0uHm0R6pkzZEU62CMLNT1r4C3X7OftAbo/D7ooGYN
gMrRRTqnE5V3+kuANKbFByjdQAZPY9ffB7tQeAWU/nB9S7CsjunpVkVUwdviCfelutbuGcGUxU/o
aoCYgKKxcVo6eQvhiclsAqOWUlCEHYsoAsUpeDbhHVIpcwu7y5p8QyalHM57YrgM15kso17C2YMW
9rSxL7W7c7mxYTD8qeze0f+7nADsnL3MpJoFjMCqSdU3X0vVQP1QpkUpZtE6LbAASs5By8OH5FQL
ILTbUk5KVPvfRqCgc8WVtp5IjymflZxymS2OqZz29oH3xVipbHZmd7ydqGDZKhJIZpFZy5AftswA
8b1fMZbbg8YFabzEwziNj7B3YSRjbGevMQFpTMr09PQIBpwQfbCKyhNUhgmyT8CiSKRu5EVyIaEh
gNrtw4VhDorrp+HV0dVa6ta7eMNan0SMMg2rn3n0NA2ABZMmgzxORFANL7YH20uKv3t/YnfhshTw
Fsb3MWwqN0TTlMXfYmMbc6gefkgwRfE6o2exc9E0YwQIEoQeqVybBd7ki5vmTxEREZSB44UPWneY
g5aiC94qML3JsEPZdJXfdH0wG1WdgodFawxQgkGBKQ2hOWSmMEN1rjyMUbRpPRArRfyOjDNur9Ha
Cso1kulABmVavQFtW9DQukMnRGOKwvucVBfvSdRlrz2YHWnZaI/q7Pfu1558/MoHkferb9QuzvRw
7PPvflCMU6WM3UZrc1/0RhP+P5W+ipdjRP9hMHZqDSXnHy1+CpwgaNGVdOIiLdrjTOyT8xJFjUuc
p2HkYhcpeIrOniKSoBfIeJZF1nsT3MxUC6dPvpXYnQt/0SvP0MmLaAzoy+LPlezng3bdhUN6+3jx
0EAlYLUSaX/Kvq8g1r1FC3bxvhp3R0FR28fzqt7vJ2fB0ydK4Z3lSJVbUd3qnNjf2Y0uMX3nijQQ
o4TTKbwkhgo3CDkNs6NtdjPhb2pgE8HN6hkff8com1gBg9UUADB+hEdoPg8PZXtrSPArY714izn3
IMllykaCwnuCngadL3JoQXApPFo53K4Xs+uM8kI+SdGRUZhC6Qs3FgqKHdvm1zLwZhDOq2d1auhz
krG1lvspfndN38Ym9hXrAWnyYdysEutwtTa5Us15NSI5MGmLdfGplePLkgw12RfeagxO6tRJY9i7
960IXPvy8QYwCm5vl2YTa9y28eBAO3k24F23tvrOSB4qjllIT91nC4IaOnQCL4mDA0TYgewuGJtC
gGTZ6NU28PeLtcid69qPu5hb06c2XMeg3wEHSCvmJs5kPLcy00FLhIPYGAZGNFcDAFzamWck9OcB
7B9FMUeJHz6qcf9WDh/H1p2m8hX3V2v8hppFBZN1Cr9LKSBUoiCwvzIF2s+x8lxhltAC+Qc/EsZ3
ETEi1wUX5SQCmhQo2n1WjzEsR6cMpMEqxWnJ4ihTQqJe+31GWFFy5mo/6tubR6MLNVmTqrjXTBJi
F/YqmXlfK43XXwFlP2LBX7+8BPfkm9MJU1SqSY7uWoGPsjhSugyRs5ulhSPQm5xd/nuRYyJ+lr+R
/cinl6Sv5fGE6pQL0IQz4zUhS0X/bbUGpQJJTeS6aKLDT8X+/JeHmmdl3pzzE6sGhiq+HFpxd9Ji
3+t0ls8JHJWmxfTTPCq9WrIqlStTDYyMS6D+9KMxz+OGFRfey0pcENNBsI2/OL0b3xdD2iPIWKk3
YZQeAwHKoHYSH7wluiwRa/G7/FXTiJnPeLWeOs15oX51/mNHAoeq8WResCq/S8DlSWaboeucY2lf
VaIhWM88HxJwFO2MvywmnAMvNy39qWUw0NwgLVU++XPaDOvzYcLCCfA8iuzDGD01hToWcBv/wI9+
pRyXwfJgG9DA4OAtK1yVnJsIoc+VOKB8Oz+y98Cifk8vt24SmreKIiy6U+3kdTP59ALYw+0PVV23
VZ9u/Um6i/lSl4iNzUJ6chHPYe0TYyJ1P86gIynMt0aMCDAcrHMRlyAEzCaLofNsdo/4GcSUzF2t
izJRA/HxcGNHv9/nfIRfgib8IYM7GZ3lZOdbUItiz8WHP49MqF4Dw/GO4uU7w2gFwq2+HchoUcSm
FBdXAcNzF3OfqPLysRhduRycqfMRNi/yv3LqMNhfhccmvT5V58I8UfEkQsaVUndylQk7NeY8SKpP
ZGIXwnPONq1lX5ANUy3gZeTnoquoEBV/dewQbKAG3QsRGRNxmXUl3NeL3TD6+dClcltw0WJ65Df6
U+JnwtumX3zw5IhaDg9HcSUjgbshKmXfU1W/oLaE6gaRxCnazdoFvSn+BIrk1LiAyHC33kl9ntZA
kqjSG1h37HVez3eiEHUjqjDU/mUaWYCT9//64999l+VtAIIb0y8b/+so4OcKuINzwLCW2H//NRLy
poc4VOHmTDP/j+7fZnjEBYNR7Hna96chKP/LNHL5wagD0oEvgkmsDHWYUnJ9BLIahPEy6lPwylMW
HHtZeoEN+JlBNBsn0K7C+Dtgq6oCGmeOA60SGM179HwdRuVfPLm6Xzlsk4eRVuF3VPNYtfgaLME/
zcetSxIXJDZ9/PABOv/TkbqEBrPr2snL6ExLine1/EOgTAT8wKFdqHI2dZppNAV9m54AYo0UfsLt
WPYaUQdpvOoVo51ZctYF+QRv/Sm3k8viZ1EJewYBnII0A8e38DVGoeUfzKvdEsZmGfo9lBai+hbe
R9EeLIAUZkg+XQm0I3feTxvV944hFhCwV9xwX6K6xpEsL8RUvlL5LDpnD0DbBhVbJUR03Gn4uv+o
206XAKo+w4H/UjzaAFrxrf/1fCpPPm6/udiK/v8WBQ4dHD0nYwr54alvFXI0taGQnN3vpxZgiMyG
/D/Tlk9OplE2omA/ogvn3V/Gif6JN9mmriLecELS45hzayrWmpw3WWwzhvC+7YkRXEd4Xmdqz7bD
MsHKQUnxEh4wQxriDVvz+eRTZSdp+jP6lJVp0TfUo/iG8FhMkPFDdQD2PbEpeqg5uM9qbTbeDFKi
WHSr7jWsVS+9eGtyhZA+LZpzNYSWXsKYewkUol0HP0dXEWBxLFRQJB5Oc/eZDkxSSvpu9zqWrwos
FtydwQK/dHtb5C+531hZUOZm8HXyDJR08v5h6zquL1b6gNCGuHWtXCbD4fwT1kONrr65zozx+FT8
qDmeauQRk3kwsRxh/kMqcUst4bTEZ1Hnh6y93/WCkQTZ9xqt1VVOxQbuWpsYlDZUW7clqvcWd0cq
ANLsfd+1vHjlXrlhPj5CyHLbksC25jWEwKntvW7UJftCDHIHmabb+6JTdic4CFJxBNMbAAEn80E4
pWshcifraxmNKG+LRPq8ntPJSJjGldLRKb6/VpbgVttENn5rniUb4YluydqlgTR82ufdF7eSeYcK
O/RDqGSzlmTOZ0rTR+tT11+nHjGRdXjeoznpLYnULJMhLABInnqooY3wsVO71IjerLRmJs8TRVr/
dqZoUo7nqfbSqWorKNAaLS30KqvRXlDWKNf3XtNUABapbCOwd+Uoq9VocI3UZ3sTiJH/P2P/DKdX
ClQHinV0DR4p9XYUxvDRsYnTTIKfZ6Y6r5PlBCuxekQi48f6wrEKPXlGpFwKRk3GKksY6RlIXh1J
r9OMjncGdO83xf0P0JLFrQBxhnQRYv9djDKOXolzMJM/nOHavVTOXhf6D5Ep1MIW4QPGRK1IqLg7
P+3tl/CwjLZElQQaoRp3vz7tN85h6xwD+6vvjqSYH0xZu3Ho1Bt2au3R4PxoeOD6VEj/0cX5vAsS
AcXdhrAW57PQ/WZooIxmKZJHq1Uy+iJ70uAzw2RDj9HH9/BKW4lFDDLbZb0z5NXlQOsM2mo0vhlc
d90rwq5Q1P3NMwz+UjzwUv3Cg5T5inEMvbRGT0hl/ZARcN8j0Bm8Hgdo8KlZULeAQqdfXo/vKm5Y
7IsHFBEtkT18WhMts5/9G2leQA1dsOFqo59aYJiddlSjQ5LE96vhgv2mT0zEOzDEcqm9ExOiKRfj
cvHoLlCwKRftZakcqqGsWqYf52bXG8dx58m87d375qSutYP7b70e6F4IFECSfug+nJPvdJnVw+uD
2+13sJqIddSigimmMD4NU+LjakoH6vUGaa2owip3bks0fDcMB+hpcWp+3wS3XebS4dl8RgHye1Cv
fx9qMmtXUPf152EQughr0J9Erl9RLnh4QIjVejoDca7snWAZdV6lpEhoESqrwbdvdVlV61EZEo8m
D/dAyzW0ARlBiBmFFAqaUKaan5haQJylh4rUqFtao8+OSbRO8COjYIvTEQwyD15o9xPxREy0U8dj
l3J1a8Jcqau8PmRUZIFpYjE/0iU+oHCAlIwlIYuXay9H/CKTgBgrIsuVlUK5d6uj+12f1cEEylKN
eKWYKWgMqLylRlqrvmR6ahS5cNnYXQzktoPZRNi65RMlpLzbStLS4ylG+A5IJN3hZKoAfNXBJzB1
W8OWWBgyafHo/PrCgcP11YIYd9onJzcyyE8pUJx5+FEK7A9+dyg2TKBwM1slBmdMLfU2J50Polpe
1HULv7z2in/MluKGHE+le+IOhXgLlnRFiPLb6vkGbKPYBM4bSIiy8NHkMaKqzg52lZ5A4B/ie48y
a7S5+U+ZUxlQ0+ca+kdgOfPEIDqfIxtOadPL37y4CVXiFvY0sKhKiUkHf0InKzu6rs8qy9+hSsWn
ON1U8bcY+egZouJIFcyLgRiBlv/kHUxMD+N5wPK/FbXtGiXd4X/CPGIYanyB1ErKdXG3VnfcI5Ow
XwQ0RfZpIvjJZ6ZI9UUGFuWcoqIkoiB6xnm4fhH99ZC6k/65f+8Mx3EUX7iv5BRi3vWxwjKIDjLf
XN43fTbdPOHkekyHC4fpJ8DrLNkblNuLUyNykUvEvJXWt3UBv5JOvsgsdd1Drvwq0oHgDBNpaXpW
3Y4VACwNmwU7/P+wj/ShGT2AoTrZs4rMrJkN90jPuSIY2PuwVJ2xhpU46jZoBwmSdusE+H/CemdW
GkEBS0IC837wiI9texN7sCASd+n7wLq1LU6OT7I1jTNBjThncU+Ou/LoLf9Kkg6J4dn67pgIH4qV
uthaK/5eHgymVaXd4coTwBQ1vMcrBOFKBfM9BYwIAWHaa4WPmyKTJMhRvRxQ3kbWcG0oLs217xBy
1xjrxZ0Fou7X9kpqQQxy8UfcKLjhpj8E777x+pgrds8QXzK/yxMBnoM86VN0JrLMn+Qqu8bAkmpR
SJF4GsmvN0b/2J0y3kuX9iaoAr6ERGwnc69PpUS+EtW9MiuT2GBgmFZwM2+iH0z5bm37K1DbnUvR
eWFivFQmqyuYfWFnm1hUYQBaNVFQ5qQV/m4/yJ/wIICag7jzzoNFWoNuCsUwiHODmxDQJyjDH2SV
UDVv5kVDmUlDM4QJU7E9BOIb9QZEpYRtOLxM1KqoEBaNkKmqcj6Yup4eZY45l6K7QXk1xqJpABGR
w5EBBmpqjJdEKRHxV7Ut6KMRurOj/KJH6SdMQijHAu3z1obv8aDUZowDwPYYtG2UbR17v2AsQRSW
mr9Wcduhxm8+ZGAGar+I9x7319/Mq1zugE1tuMit9GaqxtwXcDvr5SZcz+5PsZbnEpSJvTzoixXR
pWWuNZ/XkgqLr/1MY9FjtEZD1jj4Cbr8w2KX7tr7Ls7fiJT3ph9YonKpghJaOm4oBoTgKZKzcuI+
30JhCoX70a643le8DslUgkLPfk/0780G0hZQSwsXvwwkPLRJ8s68eIIzruy3vcOylVaAMCowB2qX
iCpx7+XRgnUhAeA70X7p1pAIENitEO64VXRK94J+R6NE2N6MRQGtx56k8qLBTo1+tvsm0zo/a970
IRWsfuR1pzX/Isl2sSmw7tGFkMhzj5TGntHYduS19nrJonJn2AD+y+OPpeXyO9+05rP8xV/gIRHs
HTvdputTiDnGMc0WOQU1o/aHB/0a3U0aB76B2lAvf3tjVhyr8jK80pkiajyGIgv6I0+tOKQDrdFd
v60Arajy3yU4kfEoZZAKWksRZvFgG4wsV60Qxpo7tTJKqGL6Aem3RrFU9/3WSoWJFKroBthZU9nl
cKcIoNPT8c+LmyvwlKHU3w9f2vzOSllTLRehAiQGX/ScM3+x7QwzFDT5k558RWuMOB/1HxboNKGf
PzfvgQw1FJs9X6Q+8ZA8MUx1Miwb8rm1VFRda5juLnjrzfJte72eQRJicNZXWa50FLt7tWZEVFqQ
xYlxNBScfhC8YUV8qUkFPHloGMg/cWrqi5qnF3Y+LckxO8S5D113Xb2DvAgjPQryoNYTW7XTi/ax
WKot0LzlbZ7EbcBTrkxLbSSYVUzSmuf/n2S3ilxWaKBQjQVAK2geeJEIHe2zWC0PIwpSn+NYV4mj
mbgPeFr2a4h6XdwVaTZwuyQce+qeESD0+cqVQe/LfGi934Wi7DviDkUs5X5J8Aq8B5lb8iMGU/2a
U7Cnxz+MwekfKTRiHDK+o7O6RbXqPCfcuoMe2MLSCVJ758rDCatB+SBXv/ig9XHd/WSBunlZGBvn
SIoTKk0rspCrdMVBkmaz1bxWtBSuI8Bz9iN3d/+EE9/bYDqKTzbO4LhNejYJCRVr9iKCHOYzNHW6
ZX6oY92dWrsUtgakdwH229cXUGWkTWfJzLopHF5dE/hQ+FfsO/r2XQd8entOt7opO6d4BMJfNMd6
WhTl3BzCH7CcmHtkBO17DmkDJygVY89joy/kUbZmLDCXD/1KGbGJVRK9uTN9KrjsokDINA35Gdop
1MBqzyRgZRDh7r0ovlhBOySG+vrOgoIKDZZBYNOHZIXeNa5frsEprVRpdKcpgCPH51b+Gzm3czEd
REaw3hTQYo/g+cNhmHRt4E+oLp1LgrOiGfO2jagHoSmMfoY2JUJW0NvjxLFIlWQd+duFZjaiIpbD
L59c5c9axpbczY9Zbr1UEj5FQ8qinLF9hErj6vTgOfEFTVnpdcUpgplwG20jMTfsxFYWbW+KqGmO
EwyRe72zfzbaRQMJIP8+OmmQpYHN0X/TAaLUGaD+NWTmcoUXgqFVY+iqEiyX2KildAsjYX7nXvSo
0jdYvtg+NQnrcPYyFcGchjs4QOLd348PsWxBsqyE1FbwfbEauVXR/lZAXAuuisKnaf2iS1DxEuJ2
OHd1XO77KNqlrVPQmBdQ57xK/EsLwvea/dHMz1cSweFreeSp/3ESigbMXfdH7CrkV31ZKE5xJ4mx
Xy37XfsbPKe4Zdi6T6W8Zd9N0P4SKknB0eLceus42DgEGy8EzeKlewEz9mVhQ7LXekpItQUSDk1t
866CZP1c7uLlSEv/vRtEmqkF+bk3Xu2Yr5Pvp2XfZwY/GWb+VptliMkfulpMudjaFDq9R5+MKjLl
9cTW8lgEUmYmXDsIweKPhh0K1UrxjZzxG/Iue1Z1aWOSSjL0EsxtYaLuXGJnwQAd+NVRW282fFdk
K9z/jhM2rDct6JDW9Zg5ilH+hIlKeh9ANrFcQLmEEAdffDOroxMuENg5Z/U5MpE+V/RQLcaTQ/9R
wuQS9U3xeZ9zJ1pCOsMYar4SGBfxw5ehpftyIs4zH7u5lJqIJ9euGhFXROj1pAKMmlZ+bu4OKxNE
ANw5tx4vn1YpoE00QcfByXiIwxd39+0IaT0j5Y82vaBGGCh8cel4XeRRgY8BbJ8y0rxNZdJ4Jumk
PGdlH9FmMkookFxVDP7LRI1HlIApf2F2c19oYfo45eE6LHadLU9+GSrfTzOrz/q/1E9CDJWQGIri
56Oe5SFkLLyE5365GZYqN52vfxVFfEUQXsUljj+NFZBkivU2AgV+6yDG+tAJHirmBIobkDtrwEkX
pHAP18QrI2NtwhJFAJAWxKvXrxweP9i3L0R0XigS60qrj2zgypdA3lrHLIceG2/jfdN8L0hLi1zG
INR6pI8C34VD1SUzi0LAyfmceELX5/x1rGKelLVBe5FWhrUG9LPH8c9B6Es8e+cb0gznmb2gop6G
KDPdeLOH16XqyktyFAaiigE+sIemJvRFPmiDpqd/qaxfyM5dmBjrYHrt7wXnI17dZDIK4z0FP+EH
G/gyeQNIPRqmTyVaqI1oy/k+i5EecSN7iK4bU+XWAaFMnR2w/bTRAAT6Rd/aZa2wx4QnheqZ11E/
z3EpGCgXTczQoW0f6LVSooF0pv5B9VScLS+YsEb/09iA4IkAWpYIQbDYFFovOinXj3BUnxelINE3
xEPimmGwqEmc5tD3dNeud2WSb7ssR2NHoIdeZq+hGGEX/gs62udButBw9Z231F4LiGvdstsr9a/m
6jZok1YJGJAGqfuGEXX2A+BeREew0mEGUBJ2HHbMOsNXzF1Z1JAOhaOShmsU5DPAP89Hz4vCJpI8
GiAyjT3KYjGHcW95OsD6iu0cuPlWNDVn8iuBBVS/DYHchY02YNBBD02pUxMHLF8alXW2WjpK9qQr
Jux6oB9HHoYHMu8HGnoVeyT6/kYqcD8wdtiGoXDIfPB8m95FlQBG1C1Z4oX4mNKRXY1DOeXoFwp6
2Ud7iFbr/UaJrwp6PS5GDLbujN8XN6yGkenW7SLPJEruAaS9hYhOM/UwK+29Odtc+aPE4T6lvfrt
lDQSIbVeCSiZ//fCiYzmKcIJEh+ttU4sH2DBYyWTsfrrgsaJ0e5Vr8GcvG2tcl+uSzihZA0qaP56
bVNU2qaCehJ7KURbj/2d3eyRVrX6sEqPJCuTg9WRfecZTwkq3pPniU3IlsoNDsDRQOxnlSLUIQsK
UD7urc461ETRX5cWHyuleJ5x2S/jOUVdmSJZJWFnSdADPViJTp5DF/g0WjbMA5D975fcSoFZxh+n
Cm437SkLuWwfHmm3lVdfPgy24LUv2cdJmgVlU+o/bCcG6/86t3CyAyF33277dSDWFQnU6GWC/qqG
m0/9vRKEOkrsR2e/qAONgm22xfPFJEfhT5WUQ4cnMxIEnhhN6soeSZv1F12DQJP4LoTz1e1lIry3
bsxZD3yDZvOlbz8XLAWRhjtrJlokcvAnq/EVSWcObCETrxQewaVwsqGFXlZeCj1zuQRqv5MaRlGB
igPVMpoYjnT32XFG+5PJZXsJqLglMwpur+tVIqf5pywOA1xp7PB8BmNUREbejhV3OXjc108NmkxT
KZtLm6fpKkkoT7e4M6xaF2L1JU4bSf2tk34rN/mZjq3kq749PEEOMRNpJCf7WWDuRM9HopKQDBSS
rS6J0Ikak/QhER4ndE943d83+ATONnpoZJxXQrRNgl/3lQjYpfY4XFgRF1MiWuI1a2hXCrOOEUzp
o8l+Xib/0DZJaU6ljckOLajmlxaDO2g0Hju/okcvXGE7er0hSoXay/RfHmYYkKSNaNgoi0jmuOb0
Gua1113dh4KDVodwUMSO7ZWaLpepPV2MeklOMKQ9P6g2gn4IfRyJAIC7W1lCPipbRxLAG4hf8gPC
2O8Mv3a5Xadk/5hl1k6omEJ1ahyNoDbVqLlUSEky/79Ins4PkRxxxigIlmqlMvzSY7nPIdwFQt4j
UHYkWAPPrNNrO6jInJ0L63cTrEg8Jr7hVfx3A8zx8tEV00fBhc7VnJ2/JcpU6Fj/txDrnQMnzwiA
gTwSbiHcF+hcqLKbYF/NLdDfn2nJlhbmgBQjlYFBS3hdXnYZO7BQdHMCRRR0jl+70QyzlPjmnhk/
4uqKcUHUFaipqIzM54zj/cjslJRtvB8UVpPuO+yHhbXX3nq56zGhtsdpQolPxJkp9U34Bt/edK+V
Ng8MA+FkzOwXRSbfUKCxT4wR9sWPVUPddZNIgmhhy+RMR5nR3R5hy9JZ0di7XLq1AhRUu+l7PMFc
V+JSqOne6LYolbzx1KkhjZul8qdT4vE6JJHwDQwGCvxHSQV0U7fL9QtMLrf83ZEepYEyKJGsUl1+
Yghgz0O3czw3h5Jt3hJ+DxckJkfclnWFD59STc3S7dYPKUApyJMLW4eO6Ip8r4elWf/7CKdZW+nB
iPEqhQDk2lN+kgpu9Lwu5+7YBst4+TcG+BHmSsRB47x3nagooLQWhDfqMON9ZzFZSPkeM3ImHvTv
GNVME7fo3Gjh+W6PSUaJDrU1DwCLtTcRX2rJ114HjT+trIvXvIuSGU09ihaA2xcUb1s7r8BC24zr
uVLCHOqIi3KRPYwJfnIZBXpCPWLmfUw7/yNN+D+rGtANIoAct3Ty4nfItOfieUu1+I/lk7msqPrL
+zZLQODhFUysqaw2jOGXN5JzljCaIH+8TcmCuA39K7qwkWCgpOcIeXE5zzbt0rmlu0dUaJArcNML
MfrI+zMyUd80NBLD/oQ9sSRB6cD5+iVVm1RTWOLF6rJu+g/7w8tXEdFJFDlH37CyWjEnEvRuPgwS
A9vMCcT2wE0N4wzfc4gCGkOVy9HvzHe/pStGmmR5yTfTb23zMqoFQuneCyJaxIhpAvVkKcpmaWcz
5YH5cUqz5luxnpSxDcseCvzsh82rUvjCMfG8CoFtr/RpUS3OETjiB39pawZ9C0Rt1ss+4RZvbgA1
FEXTAuaEaV1tqyyJ91cBopr5OZs4zSuB2TJEV55+eyms7vwBDFqgXeC6H8XHZcYwXpi/V+Aft1wB
Unt+iIHuTSf+GAHT1nVk0Oyo7Pe8BLr2Vj+l0qJnFkI0kkQlBdebHzXlGOYI+c5cdqCMytcr9N1z
1DumocSIgf7mVuC/syNUgafe1gnuU/8vIL+oKfa/x1MWjdjZhUxrrjFfTmI7QPt7k1fXI/hobQTM
ZhW7cL1EJdT3ZVS1/0tfzImRlRdXUF/FOowlEnvy3ZlCq8+Z5UxQ6+w5aGrHq4XrXpfS3tF5XtjC
7X52XG+vQ9PdM0iQ0wWvbHJAEa822/o7U1H8jey9IAn0OamcR8LNUARYqhA/pzzoYgzKFlBOx4sM
iGT9AoPGy+Vk6wiwbSJAJi31CnbO6FXbtaLJ88y+iKMcK4B9cw42GJsA1kDg9VB1m2Io/7J3pvgO
DAbMYXcBI34kP2oTQZ1AyU7ZV0dlK/mMEBg9OADyKZBzxwfU+Sb1EQNbqUwwOl3x2YInn4fvPJ7M
B68WwuVh9s2Aq9d8yN+HApK9YLuGZLH5HwFhAD04cqQj5SA2BED/xPfRwWekC39dSGr1AY7xLUw5
E8O6sdbtGodkiHzno5KcubpWETxKP2KaUiEKc6543Dqy+n8m3oEouAZuL8su42JJLql/eyMqNmdY
o8EARh1DiW5Umh/gINZ/wiRVm5iR6ilRNhUpnyCYICfWSpmAL1GcPC9x7CVUY+heM4Pj8hO0PRmr
OmMR7POYeiJ0/KZ9y4J9nytDnOIQrog2GCsSMxgY0GnQoOdFNE3suRPh1ARhTIj19ppLQly6MMlu
r3Ke+3KwHCQ9IJFs7pBZXQHnGAyNe/OuVYly9lPHED53ztQHdRJ6NIouk95OAPc5oAi4Z7wjkiLL
01FC+bQzK7YmaAdLmbvi0i7AXS5K9egiNMXDukiKiqmWdkKNdQ8VLdXxGvmWLASH83cmJ+8Qbww0
SE6kV/QvPfACscAf302HsTIOnP+B7OgQxmpygCee19y4pYOp463MQmTXnluXzuspo8rK3X+MZuRx
3ICY2Z5W7sEtUqBDPKzbRulsj/tWY6xTnboqtVMaF2vHZtT2c+nb7CbOf3D4c075buZ3HXuV4M0+
T2d6T/MTTKuDlU96kgPlqfa748kocDS6qBu1UmfAS68E31xoUw5NJfQLD/XJPSwtcgC7lF4c2CiJ
VHTc7yJwBpvao2Zk8OnDOw8pHTibM34Dz8GL6b8C9hLlTYB+3X/ZZTNS/HFU07R2VHbmWUquET4i
GraBnhNtXnKeNKtrP6ndCw4NA39ra29wyybkB5BSY3/P8Cpb0ViKe4eqLGF9Ip1AyiTX4nP6eI78
RYBglTVV0lVtPJduHA7H13ed5chAhfNm8OZxbCcKJqtYHWm8JpBVxiBoZLVZ+C8CQ/nlrRw0fITG
6WGW6eVmVyEHrtGQB+bkwLteXDA2RuFFMckZckNCHJKgvs2NrEBaUOzGwGJBgCdNX2zLMguVkJaU
RyM2lO9z70l3t41l+n6lz0y9vbw/75Ic4P29DmKSU/Yi46gG2z+ZyUJnbm4kzugyIA0eqWx1wuES
TkUcCEGDmEZBXV4FoOzw5dgU8nda9ExjmKcfRXQQ1SR/iBQ9HhI3vr2RYcTB/Im08TzzOI803hl6
UlqIQqUDwALwoZsg9d+EkhuhtSgjJa8DHHMgXr0RP7RxRUhj7yR3w1W3cMV7/l3XtJIB4xjua8hP
8/+tCnS67YbRfrrguVAqEHbCrn4EzL6zYNpY98MJ6HaUw14jGatur8whFxWie0plSutwAqwbstgW
aAgfDd2Nmzwwq59LDHmj6UnaCzz5bXUqD1DWsmQeAU1maq4SpcFLhD+xtL9qZK0xV9tw2sCGySx6
iC2q/9XRjVTef/HtwlmYbwSLkLBW3VZM0D+ajaV3IG3t397lXtw8meXe3ahetgJ3kMabLAVMxw4M
KK/IQhK12mY/lKBi6phmz9BkAFY9IfK+QWsiGC0nAxl1iIEH28uDJvZuUepC/AYIvIpbr9PBVYVQ
yWhz+/j9ilfdYWLgKnJvXe2ZFzcSG4odvk+G0w+2MsowvLjPeGC4Z3hwyyV5Tkni+ENTHVzdMo7a
ggLK4qamZ8XPgPk/TkCAk7PM6grFk9JR+feFdwRe/EZWXLqd064OsMv7mpKXnreIBYcPcyyeCmO3
biqOqtJ1cgXYx21coUq1R7qCd8BHU4evE6Sw1FlSEfv9KOmnb8ACES/XuMUnCwt4FUPDsU2zFKy0
KsuSm9t5X9HR+zm89Ic0yvl/pR1CyinYkla9oicW0DLeop/fj8nKM6GAXds0w4n7SmS+JByIUiST
FVATLFZchRiuo8euxv8vXbBdohbHm0AxyI6keVrzvW9U5jGyesx/UWFXpG0ZBszDhC34u7j6DCJa
x1S/G2Fa9NvCCdBXg/6CeLl+kIJ1wXrRohQdY8Ub7gxq3vc7fj0ZgxHBrwfmBqZNqX/iF15xiLpe
aakuOU7xfI1yNwN0lnU4Bie0XS0S/+1Oovv04oYjPvbdTAGIuYwvS8zqfEMATvgoh6Pjtpm2SkpO
C8GcEa1++fAyGcvyy68wWs0ba63OuVG1ftIeqiDmryZr1Zo2RdBcy0MD0WvAxUYdzM/RjN41J8ZN
7ZR8zD1lyuxjd01E7tuC6cJwSH/M54WBvU7IQ41o3vtK+eH0QvEWuvEZTwILSpnxg4BXixfybO51
5WkVLlCOKvUfy5egtQ88HeSX0zd421QMsltqQnbU7seGTfvPOGVAGfE1rXfAFc7I7rlUfNv+GiID
p9srsWsi4CzZ/3p9VTaH5oNaUTQo+Q+VkGAzyU6kWyoSW96Rrz8h0Vsk0Gy5J1742G2CN/OzDekD
VqsOp9Emx6d+3aZgCov/EGNtOU7GnQMiiqE5KYXURnfNvhNuTAvxQyOgDxuaGa12UVNMHKEaZ+UP
YI4iBlclD/cu0oIButOL9mzqz1yOfIt7IRXGZ0OV1rUS3Gni3Tn6buBJ/tSm3l6I9LZKchohjXEZ
7jb2cYgQLGND/p+kr2Emyqoq6qEcmEk0YSZA3/VOuHi88aPjH2VDo/JOy2zU010xdGs6SxXz+HoT
sHhRUTBmR2OsG3StqBB5/d/G4d1MAocQdlzduKj/574KdxRZ3gUbob75eaBoJyPAE2x0LxUo8X3p
QFAoJp8KCCFHPM7QX1v9wczZnNOmyifvXzw6legAUeYyIYbKEgrGR2siCpTlcObOugCZ1x+j50+9
R37tmAYSLNjUW5SxpGGNqn9OxrWac1/sX0E6oXmylxF4oO0CCtRWgIhof89y/CQIqONM4LD3oBl3
VJxyMtzInq7SWVcHpl8bgdfICvNHLkUUuiscRZ6b2UXP/+ec3J3dhWr3txbjgRxm6lMtvNSBrJDd
FN9J0wgnq3CyGHXACwSOEAOPU8zZTQOO2+6ao7bi1EaFg0R85vBmbXDtGVOTx6gLfCrYYCZ8DfqJ
2n1Z1DD3uREL+d2KjGt/cclb2BTBfaq+Lh6iMk+Azdx5IycnT13gZwHknJpoU7TsLOV7UH4uUK6s
RRSbcdC9clQyop3iXEsnJgZQoPAZeIUU9dFEqnCOkIAgPkH7spiJcGElmAtj4uT8tVWVsKW93OES
0LaiNUrQwkkSonrgv088r6MYCs4F3zlAklCEBky4M/psWxG6M+YF72o0O93UXDDLYKW35PXnhoVx
k/hEC2yGFbwAcvzn1rk+c+5ZbKfmfYUyVOOiiQYhWnif2s+3RW6P7OawdRRG1eSaK6A8JyOW922N
4vS36JG4gwcMneeLg1hWRNJ4YXbPBHHkPyinFjnL2t33AbWafJ/aNt6JKXAZ3QqiDB4M80DyN2t0
1+IxOpz4LWaTS05e3jgA0ypclhEzXB+koeW5IxdLO0dso6A8+r8xCrTLtXFNUCrwlI3xz5/QBVn/
kvAsgJt++NqnC5ms2u+CwARfLVIQmobXG28whQLR17qkrsedaBIyi4jZXJP+yEUe7L4bB8GbfFQW
4ZQoepxYQi3j3rWlLCLinJ8opOCsqPNh/jVFHvzskqCX1G17/d1uarpaubIecwwHQRdW44qqLhI2
8yLiD7SDRarPWlK8SzUjweLoLn0IYssMPlem5X5rVmScQJ9fo7G4p0YP+RVOQpC3kgw/oX7hKnVo
w0kd6RwJdGIXVKJZv2azMILkCDpp1n/Dh6Kxsa8G7bZ6D14lTIVwP1qp3YDuFnDHGTNVTxkUQUoa
ytcuqtnMflLCsvO05YP2umB1zSyreOvVJGhpamXYP8PiqL55ONBU8okvHacCs3zjta3CbtXqh+g9
mQTEqc61uKgCU6F3emlCOpPNlYGzmT7eejHxrCxasG42Pr9+Aap41hEL8GgjciKpoznTZm1MSqIH
8dcVtsz5mTwubNUoGYPMdGSf9oMfDMWlJ1eAUVXxvpBfpon0DIXMT7oyXME40Y/VmW12C1kgrJsM
6bWGxQJWd5/BYBHS8OmWfsJHki2LIpANBRkzHyNFroe/lkW7a197ETTDQVV1flwA9kRAlGshTu8u
JFX0LHY2x9PjgpURo1keXPSzTIqSuKyfvGMc8Apm3dEHR32mE2v42h/jiAKQ9raIu7ogNej0sGqs
vO8++yT/agWuWZoyEAWULIzjzAbWAfQ1ABf4Mg3hunSYwWXoHkmFVPitYuYUyn8d6jHbsz/Z16hf
unlsY+iyG7sgkxIO3zKVP92L6B0kbWfB/eBiAQjGjGZS2XA8PRXe9FSM/VVviEVpG4KnFWXcUDPA
AXcjjFJ+pAK6ic+xntxYjWhOWjB6SbxYQAXcczUKVoodD9UkrB7tt3MYg4QIVg9XFIQd/86ZaC7S
ibDhLAbBqxTFCe7UehwmV21Bqq8Tb4vqSVeQG0JqbxfVrt1nhaQoY4WsA+of3AICNKxsVE9PhA5L
8mTGK/IccUAZ7U+DqtLThij03/A1Xr7MwE8c6YJVKX9UN6UMq4Q+3RL+9Hv19vxYSijkgbb/PmbV
0FMPZf7wwkYQq4AUSkXpO27inJHor166fclz+8FWzXk1hcjAFNgQIg6CUcQRtDpqBWaM3IrRWwud
CEiWXStW1Pa5jHK8ULgJAq8RCCesgORl53fUcJn4yxP53UVA/iDZMuRvXgcf4X+I6IJLQV8/ysr+
QVDQFn4G730IcGdeTvD+1hUlYw+WiHRCqInvxL0C4zyLLWTiJ/ATHa7XLk9XSFAfV+7k5DkAnXgU
Kb6Pz3OpD7hLvADrOhbfbF/bcyfjypEumX9Kotg6ts3Gwf72T21kU3Wr0ITikKMwkykVmj58wBSA
hsIXhJND6zdfb5qukCwahrjczbJ33oQ4EOj6yRZTZ3N5M8lG2DLQGN0xxGM3zf1OWEJvyjyvVOXw
F1THQZvEpfAki6Alw99m13CewG/vBoTqKF6Cx4k1x+WcOQSNEfiIaRT+Th3TR2V0RkMxoZqKa1dO
Tpn2lleo4X3IGER+lZVmaHclDrTfMAbjNFWTekoej0BQ3X+JRlKMWtOeTGMBQ1hQIneYzs1mky4R
0DPf8j+ybjZXQ4iDgWqIcNOtJBKwTpkURzLwq3ZPgqrbF03OUyQX4E9bVlle6QdmX5G9dbFU3fQy
uTBjVCSzweeLGvR0NO6S+LLdTYCmvLguwYO6+BEUbvb+Ffan/pir7+v2zAXBltnvoprjvwNwKDSt
dCJFEy2hOpuzxZHfl0p+0loiMamvFX0ul2iycj131nuJpXOIi8z/XnYXilKuAZ6+/+cGuaMr7yRq
f6uKzepLNLch99ye77NAXdWG3Cui56scu/CRvtmKk1kfGGEE9fqDspvs81amf1VSNi6s8FRhSdzu
19GZONW8KozbViK5GRIt7eepK/dZo1YJi0QqWHMvz/+AO0RBSQ6dSUXOQGr8Y8Gp6BhU8p8vvTZb
DLxYCykTevHRAefmzsXEk70uEWmPC6+ELQPLZV8PNDOnLNcPMSvqJwikgwJF4vHDseTBDPOTFfdm
WHSjpv4PpPxOeN9k1JQN7OgZ3CmB+NcY6VdTuNRMlQ2JCaG/SzL6XUlxgfmKrO0lhEe939jD8q9X
w0RdWZmsSvOIHRc4PwgSq0Lq7jOn9FWa7R+Keggp8DczKCWXPIwaMW9/VKSmS2EY/m5s6CQsicg8
QQfRH3OhepM3RPUo4BhsNeREHAFDTM8kLBKOa5kJ20/+l7DMMGkpjq1//m5i8+jCdTB4I9/+RbQ0
cCGb7MfPMVjhH2batvoRb8enlJ9BxLYVDnubwRxTVLLLuIvISL2jeMtoW5l/pP23aenDGXvEBaJt
gdutJIX7yXpa4uWfKANCWIWzWPrI+U87pwjFs428LOYEK2r+/QK6B4OWjHcMBwfdktzdJD2If47g
vlHf0IImQNd89UdBTZ1U7WnIgSi9hif/HrSb1dfvi/IHIGxyBvbPm19uka8bEpkyP6roNht06AV3
CkMIBkfh06EWRsYcFFEzpilrLWszRQe5F1WlMNsrgH4G9+K06N3NayNCMuSS3P8nYAkDQKynfSci
JLyGzqkWR40Q5qCqVWouNtABgs/k/K8zO5NT9sb83rzWUb1GAXgLqOTprXxOijnKI51yMmJeIco/
Mw6C65tcSoE97A+GvAxU8rtzmPxhrwy5lHma16IcN01+Hfb19uX5oJWZrEZBZxtPEqP7GXWIKTjX
e5+zZc9EbiEa7nlnu3UiqxxZ2Tlu1cZu0to/bUbZUdgjQ4urUcH7MG2Pf2BezvAt8aTFeYuhMRw4
XjGDLYlJrE27PBbYSUs/eneey0JgIO4sbGa/zlbdU03f+9N4v9AepQlT+UJnEuVsFtl/eaZdDMAg
DhjcxFWqq+sr5Zf6k4IJsoqgYbQBwwkHfNFLzqfWCCzqQEguH3ruPdKfRIg2n+ZbkIxkAU+zhMcb
1oRbL4e5CS8oJqx5cBQJWv6WqMy6tGFZ/IIBhpUjZ6R/OU7GPWD3q0xhCoB1eanKB8Ykk2+6cGYP
x8GKgKcHCw5lvAhD3f1YT0mG4iZ9aALzAk/+JSSKKrhiPqOMWvhTq9uwsLr7+f7kA3JipDYWKBIA
yUc7EbChbLIzuG77w3ahVIZmYrGzDvsZ70T26TrDo9BTipH3f+FExW60VhVHjLq9K2Fz9qHHGYKI
LuAtaqiRPUFSLQYTFkT4uC9E4T4KRE5O0QAxFH42/CEEtHhtJNx2RroZiqyme9W1avcDBLUtWIwJ
H8+3j0u05mem6ffDHhgP2HSKskiRkkmTiNSmRfRJD8Zkowp3g0QZj2uDcYYBDAZW/g1lz2pbODM/
cxEZ74yIWwdXTYRxdjkYB6zpbsYwGpYtXlxJumBUH5FB6r8xA00NZ4PsvDyDKuGObK/jS6seIu3D
RnyljDF0YwC3g+qDH3S1Cj3HJkyMQo88HKmuEJBasv+PDe3qBQQekaC2X5PQyOegQQbPNrE8yPsw
+ZorCkqmpQpeiuRTErf6Y2efS7zRwokDAWIr+GlTW+1qsQIv8JgPUt7RNjldpWYpFLQ49V9I2yXX
xP8Su5qZNtFXtoyRI9/45muPGxd1gl6shP/T5UR2gIhfWtyuq83GuRCdqBSfC0kOsSOXPwu/Y2Tv
9r8Q4+hmyyIiT/P4IUqR8X342z7z5pctl+2GG6YVUmAEoTQrmjlB5mzhFq5Rv/ngUQl/QE7ncgH5
n7Zr+otrpHq0ugNzs+j/rTtWwWyHACPhflKuT6LLh0KdbiZi8yt5DOUGlypXMW/Hrl7HEIaXuSgy
KTjc1DKlRB4zwKa/BLwVFoCNoLY5SvLFKKM9FaP7NmbNYQbUmwx5ehowjftG+9aDY8nq4rZsYOLZ
qQoz0Hy1NZnro64OR4TOmbo4YH3ZJG5jteoRCVQhIyzMuwp7ueJQzAmy+Td8r39W3rdo/RJz8yfH
dWQXfkm7V8ugW4qYcDMcb4f6Q9iUbY50innrUl7pldGay+hXg5pL0/CBaPnzJAu046fjQQg4PDiD
XXjsrOxV4JGpgaPUJToop9iVNQgYixC6LbyJPcU6Sx8SSMy7eKbRPRCGnVuXhQ1YFs455wqyp95I
vCOZo5MbI4VlWolENqAMYjhwrf0V69y8QeFxQW6g1HU0rgoer52Qxx5XKQH7+aYuqkPJbKb+IvQ1
T3VK+esSqP2PYaf66kYLeKeQ9A/b+VvfPiZWF4T8pZ44zajo+KPpjOJ9ZXHPGMQT57U/oX+cMEs4
ZhNc/rThVySotPrxrWznbcF2QRy6VAXgV6BPUobBqu57YOWOguWgpT9CRox04X/lG85e6draTOUB
nh/NnIJMuKUon/LPYAUweJFKsCk/vf82um6qHRbVBG6Jt4Chx5pmeAxJ9jCYzf5zZZEf1/gZjs5Y
SrzaijcqXzrz+ZxJnNBOA8N4lLhC+moacgvE4ZC/tZuTxtqPWwUn9zrjVNGpBYVFH/trvVyFXGLn
+FuJO8NOPnx2E1IUdkiCU3aklfgek5akpnmVCW5A0CdSVbDPCBc+Hg4YYqtxf7lQF2AdxBp+uzKk
HS0/BTpKU7xnl2yqNaHl7kSQ3xyD/SuJamDtdpV/IDGXFGF5dVUC15d6MVhnvN/nxgR2m6VUJzR/
l0xmy0UkMoSWoQNIvznn+Qgcu2RdH+a3JrhvfJEhFBIxEXJa6Kn/z22kP0ZzaklMrw4bwFXHmp0k
QiaIdLkqcgU28Hk/BMrOyBAXs8KsMILccZOyKCIUYVxiPH947nlIS1vLV7OanvEQo6fzwuEpV0HI
NGRY/qDGpL29O466A2qJKWZUCahF7wMAbSdv8l6FAzbfIt3rIjl/v+Yq1xqd7Z0q7G7pPuo+uRNX
sbmc/+MUgY5xfp6r6t7uuVGWVK4IYN/fWeeJk9FGJS1stzdtgdHoH+0zyFaJpBlyqMb9y9r3JtWQ
u78AlXdWYTEKIv4fsFWA2Sb6MgKeRcBVhxal85v4efzFzrZt8rBKG3Dk4fmQSyaR5gqxTGvwNN0L
qQ2m7rs5gmowR7CgD2UgRkIQYC/6mbGplIKBvRAFmbZZQxmoTWl0J73Eh/1f1x+4OT0LSQiWkr0T
gPDuLP74IXhImomb4G/HZDcASWYHzB6w9ZCBQrqOHwcalc2zY6G+YMgKY/jC64BoI2yZQOu3o1ay
LCYjRjSl9DEJWu3FA7LNrYx9kXGHfrMWeV7f0r6XmMugV1tZzbt9ERAqXzNDaO3eMRiS4sxxWopg
2e89eEDQx0AUcbxPQz4Cqy9LImw/ABJVgzNOijrru/95UW5LJS7J40A3nHFVW/syRG2BZTp7v4O2
9pQppkgQ7wA91oh2djMqtp57l05pOBnynqy8WkMT1z+Iy68Y4giamQTIx0w24DhhGFjGpcPi1eyP
xdtxLeWG77xh6cTysTX7kW4aTfzFx0YOW3OGXitQT5a66nBG1s8puHa4mvNFfpryvLpppxmPHJLz
UhyX4jlADCoAPEIx9/6/trcOHSto6zDHFdKb4FQMnJSLqG2aS7w4p9BLScYh9xjTgfxvw8jGSjCO
OpqmcA8SJec6LkTWOtYptLkHgoPGHRdwRh1ylJ+yPyMXRaVdk70A5RNHifB9Kbk+EvfTAb47rtEc
zYSgRBGNtrN4lgcM6GBjR9qyu8KKhymJUUUqgL1vtbLn+7+s2r6pavKcOJEMbm/sTSzfumK/tNjN
NJ6CD/RR5nw0FOz09kncWCoENVaC0FvUT+DNmqvpFliCzHcJFHNr8X1UsUpxeBooLe9KctN5icSa
7VIPpYS/0oNmwFbJgGlhOXDNhz7D6pJKQTCh73xxnLjtTN7Y3CCg6DEokcr6jVDBxNQqd+Db2xt6
D3AKCUUfrfE9mmjbxkFtDJ6SoSs0bzNLCu/M33SVJDxduoLZDO4A30H20fPwWDsA0yqcv8triL3s
6cep4IKyqWZ+rDhxjETy4hbblXo+CGz7veRelyno+6vzFcGEZGVQdpE75fVvEANmxU+Y2v9y9hPL
1Of8NozaPs8Hq0SZbmxFgkVB7lkFHViPFBglFlMVVx6ORQfIjhO77tBdRNpkf3Lj21Ezi/HxOBQx
dUG6gw9+ZNcakBf1/wAhqF1qCiMloQzHLyBg4ikzsc4P+ng/AYy6Ph+JZbCZYsbNNcC0nsevfA5a
ZHzYvjhW6niXRknfh4oua3MB2ywTM/y4+dyb03M/hRAumvkjz8aU8Sv2u5WjOO8f7klTd6mdFOf4
CfKyTv1raBxAAJSB7vsN8Ad7w/XfksrjG3Zj1D5O+IR/i2AqiNnZyH+gvH0dYWjPp/Sabge05eBf
FOdZNPjimPzXn/eyoVF8qlr9+MNHMT4xJrTKCVsVs3XXyFpgMKpXtwVr/o7FVRTZYDSLwpPvovHL
QlXtb9Ac5sMBqhDfU0caqY050lGje78FRYFbgSk1tO77UHjpsNTV3mjjaO/aQUeeKNCJxMnZ7cI+
+4+F5/LMHpf0O2kFpTDUalsw17KkZyi+LPVA4Nk8gtdB3bRBXDvvsp4YtAWRBYwW/hdL7VdBhtu9
4fUMROkQGaEIxujfBB9hTwi5p6nhyIfk2wV+pF5mYYruMo2mHI3YD7QKbFv5RTqDmT5uAnKKFXTE
6PxCMbjCSvOzwM4fn6eBkGsyWJulVMGBOUKxdu+ztToicL4tav6aXO0BExmQ1nDFz22ZcOfXJA+g
0Fz1lCfvqxNiZ1F+Ea1BsvS5vYPIH4NlrsYFCM9dxRgX8WgR8el0GZp+J3a3jyBB8FYtJEVWRdTJ
jvbSyZXrGeMLAuG+OxB4IXWn1Adiw+zTWiDYk7kdblev7RVTZhxL/LQWXsotnYNN1Aef0msCqKVu
xJD3wZuows3UCB1V+pjBGsR10MZ4+XH1i9o7Oqt+cL7BsP5iKzrDC8bW3v3zbwnsGAbN530tD94L
Bkxlx3qrO3DCGd8eJKYOjbiRJGaMAOrxtWq+9EgiXk8sMUZqPFPGrkFzbagduIKk3G1ihXI+TKwG
ipDk1m2t9V43RXP/WPCc+FkpnDT0ugjcyd0qS6wsd7ao1R916nVPcss4n9FfDcPubef2bCyR43os
F4S0YxgUJ2QuqfpCTdMCIy3vLAJWJdM0GFlh5cM+qy+N15kHZ9rHbt+fUIJlnfWvbO2fDiHLU5g+
wYVIAPlwQGbjwBfPOeBqFacsbbHjiiSZ32klMPsJqixDUsmois/jg3xIrsISJ74EAN5JN3r2Qwnx
0BuR035zvDgX6k9HY+5S9+71PDbDAjToYc9AfghgtOs1JBtadM73RRd4OAHt6TVTzSopYGKBvcv2
vtg+0TVMwrSn4x24Ijp6UTOxUIPZDuMikRhyN6LuNBVPgjH3lWRv5G9YMp3Yui6t+xFuIVN8mkcT
vLwttbQ8EidnwRO91JqiBubS4WgdFaHZ5rV6fWuXPLLV9h/VHatVQ+twNx41DzZi7udHelx4GnJ/
avrfvjPmovinAbhc3dMGIcqlOPJC9J3chxV5Q9XdYsY8vHKRzsmBAMwovPoekJK0qKo3KgwZC01R
UqWzdhv0BxL0jKzvz6yf0mrXK37xUfm9OlvmnEpYbeXvVbgsk9bpJNDurN7uZOeYldtiRVXvvJVm
LmKPxBIoWMUjWjWtvP+a6Km99MOE+tOFa3zc3kqhptmR446N3lTkfPwOIvWfmrrhQdWPmzYBgDnR
yXZE2e9YVEIZHZWSJEwVA1y51ItEo8i4M6JviuzO9uvhDoaCYvlaAsNpNA7kmPX67ULdWlbam+ao
KcVarG5Ra2nLkeit8Q8FjDIIjMG8J4nKaTWE6J0PHD2Jdtimy6hOEHYbvyeNHiADZLg6l77nJx3d
stuP/vcTYmWnU4JAceY66smY5hbqK/A4lY4sGD2uzZKGYWiXliCNEo4qRlnFkE4heqO/7oVFl4Qp
BJR5CKWW9Bd4gdRfYY8I/lUiFwup4cHUn5uPyD/829IURe6BxRT2eF6M6yM++SoppN4BYsPM/S9m
AVjBWA0ux/ltVJE5TxO81YbaT5BCcan+cWDhrptUgcuC9vpEn4ntRmf9TDvu8nQ90Gk2bC5BogJJ
AdeaDldpX2InlE6TW9uGxIM/pw6rtEKbZTtBwsJWXndqhVBI51sudhA4ZuX347sNN8ZzwAHUvzQP
PchkyknC33uRRcdrAeYlKtsVzUeZ4bPmUzkuJjVbjajEw1rKx7lVUENgscixrE3yhQbJHZ5w0GzB
MKNuGsjkGgZM4WJrEw6QuHiGPefGgNtsOqFYad+FQOmIEc2osj5yE2RnJs2EGrmRfsiP2eGRPXre
BZxIgoUMSxqpG57GayRHJxc3jxfCg0ihYOe2rl6UMvIYG9KaGt8Z/Vum7QvfNVwUQ1RoiapuR74s
tm2nQsqBsi4F4s5fpHET7vx2siDec3WaeVyxVk9+PHXLsGmoEM4+gz5Z1EjDpGRtYCNxSIvrUp3o
CMuk1NIYaCC5VFOmFkcAo8sbvTmys3HJ1aCdIFWodppesXLOcDOpQXV1qkV1vbsPqacCkzN//5J4
AC7Axy+939l84P/o1slPdsXo84SJTOPNDQ8dD3YBWcGSTrQ693Hzbn6pr3FzYW3BlRZFos3UnT6e
8a8f/7QNPI47sDS20GjWzsZI3SGTOEmbTzpSjxlmQxqN4FlU1igOx6flrLCkV0r+CGhS/Xr5ArfV
uh96jXrJMuCUx7/Gje6q5cEJErZwgiUsYXKCKcDUc7py6bqSoV0iXPybESFA8j7PbmWw4hFUo0A3
reB03N23ZCaM7wfWbyYwbeXrcZJr7LIvG6y4qRIRZDrMp1OeRsJTj0CiNk6fGHSCwK7Ns47iyL7k
ek6MfOUQ+/1kbL0IhX0Pw1aBE+nARNzH+adiPYBeGYBO36XliBbJdcmpN2XHKm18Ag/6X82wZHvP
sQyy6Z9nwHIJlWVgD+MmEGGmJYMCnniRx1a5Jb7XAz6aM0iVF1uzLA0LIo/oetmmIANEHlFZu1X1
vwG6yUlrjmBJWx3Gzxu63yU94XUa8pL7hWRBLDR7CqLE8ph8qej2WTiINkFadI52wQkWxyyU4nF6
zkE3fzDU9vp3Oxn+Fjb7JvAbEGFAROl+BWkaMMLDoIb/MxHv7+tsamFEzCXiP2YQKEpoDgTwm6Ym
Mi3A75dqeSXM4rKhtdWbVyDUXiFt7g2Xa2xsMjt4+hOjcP+5vCNSprJ4m8lUZjrphaWAz6RAdgyf
Skjf4NSaj7rrf7bc1rfiOPecD5qu6hmorKKAxapzU4fQAUfKfAgBssxFE6LvNbIFpFEJTZkHl1Z/
zVm3QmsLnUuhfmQtu1cDlV3Bx9SMycvrH+cpU3lkZ/GDR/t1qwT6aGju0cyB21ErgCeYNCcxr4dc
qZzNzkqbxJEl+sSogKoN+K4ix14PvJAyGjB0UmLzfick9rrKwbotUiN2im48zJG8A0j7uIr6GDoU
cBM6IRiZG7d22GoIzM7ebJ3WhM/gtdxvszBOhZZBHD6bxibdRPCInIbwdBDB0feOAf3UxmMHklUh
lQUuzOn3OWIJ2RHBT9CPjuOy9FFpcxutPT32GQlvUwkUP8zB50DmjdEgtfqNZjxFDIRZp7inu2S2
wx0AI6ZjxG9yYtfgJ+pTYCxMvywOlfEqIqQFjHBoBu0TiZFdhZmOri2n++dD5KDQyrkeajSrIRdC
J8ZJ1+mId+2E4uBxDPKb8V9K/74SDJAmB7jjsZn7VME4+p6EN1+Q8uxbABt2q/9imRJOe/Kp5DGR
xwctASmDE4dyHqINtwgRbVmqJ124yqOyx91HzvC9rlbbgy3YMadO9xDHAxgnjffR6dUl96bnlazP
G5hXCtPwVBVxJiCltuggTGaGLTNKVJAZTyl2cMVsHSq2BJyxrT+6InLdU+9mtLF5VDDco0F+lbFJ
xgxYZCymuLs/Fk83OoxJeVJjtU/PMCNohHh3g6erFtpCXYma1Ci0muznQEKjQ27+uYj08qfA9c17
7sAqIqXL1VUvlalFNx44VRZT6PucNRyQhBewZaJkvt65a9waKh6Du88qeoleQbhoX7+UOhZk7dUf
ZHgfHYXNcON/1+P6i3MMZhxbB/CNxXWOsNqh6GulCcbMbCGR/s4WreyjES1c69BxiV2RQ51IRdD8
Ryu8Vmz030KC73hBQV4oQdDVxO+zkUIjTlXwlBjrNN5cq79K3RcilVY/QeWTvfJnMvaRPF57lsO6
0txWPpYn+C4vChP9MnZd3NKr3OQpyImd4hjpeo8RMn+EZAsnd/FqX7jzLZnKW6rQGR9Mb2htLDK0
CMBHggRd9r+2XnusHfPlXkfUiOZCc017niMwsWzKV7jCI8SLIZEgflBO3DAc5JrWM5ghrtm9nMO4
+My/OlJ1T/HfCFx83H4xvs0CWRYgXgtTOaxcC1MO52m5jkCufP4qJCJASL84sX1pmolkz7dl7HnV
uQboefR6oNy+lilNKwbZ+/USbMaiF2a39qF2g4YZ8n6C+NrJtLbU8VVUuFpGU2tyyHKkZ2igKeoy
Zb63KXU/ofGS4WAUSuvbCt/7vftYyP+0w+gk/RVYOiRaUQiucsytukKsZ2505s1kgfExYyqsJyax
QL7hxO1FycdxxLlthF45sxNu4l1xSACId6k88i73KdnmJmCzjXOPDTwbS51r4OFEnrjwcIExhwxZ
MEC589LQyz/MVK2LJ19HLYPGd0VMu+Ie6PBO/4gvbGyOBSg3I+s5lxgRrFFvPAQzoRWlZpvkJbAS
81c6w8TASGIGsyDIlpsclzaMM7YKWaO/lmlWGjSCOd+QlNG99Mgq6cvrgbQiTKVE9smmQ8wI3SMI
35baFRSwpf2xy7Ik0JrR1MkAnOInSDzRQCTiPc0GV9dfGgxdJiqnn+gIMx+gwCbhCn05uDTFOZom
GnCheufoY8y886nqLT0Q37kvk8vxBH+N2E19SSYMslN+YF0eUTAG7o4X5Qh5WN7TYhZKD7rcUtTW
H8IOt/z6XH2KgqRPHRRtFNIJOz1nGKNEK+1/5cO/Oijz35d1I2WZi912b1NB+J19whwkWaGUErZh
I8g6UrvCEzhHDhyfoNP/K/7Aeo98n+DLI/3vL5JwTSuqwiz8rFaCPxZw6tr+X6C7os8+EhNsJASJ
le1q6oWRTtbmuWE6FO3b48OyUcxsfWUw39zaM4vqfdNCw6xWCAJ5fF3yFdFDlAyu52Kuzh/loRsj
KjYdu725BcvzJl9TaYChYt38b/SFO+3I7po1fKeSQo+hNa4W3aXKdc3+76Es0OYxHPLFeJCvlDQD
UfcdsJLfR57y18bW1rAtuhON1TdgkIcOjOb4q3gsoOiK8Th8fF69vdIzs8zgfDKOm603faZTHmL6
aV4lgX5dcDgNz+PtrGpj9tww/kHPNakK9UEJyUiO+e3SMIt7eFD/84EOHGeT3OvCSDhWREmm4aMG
80Wn8BOCbUV31h+S73dsUOKjxTR1H1YtjnHSzCkYOTqfZT9JWKYJ6u8Htyu97oLXXGxUXgtKVtkI
DXibTSlXvTWPqNo3bO7Gv8dH5ZfkwBFLb2hUdlfxV4G2hOCYvFX5Lq/QcHsKwo9eHs9eoKMWNFil
OwmGyzRvUaCJ9xq+IHv1Ld0lDKQNaetek5s6iZ3HMas9b93GMJT9eCBPnCA7L1FTnhPzPxPILWci
uyH1S7oCVXGiHiq3aUJfSOd35uCFHfkiC0wum62jkEMbb11Od+3dDs3+aDTO0ODiyNHD9ouXnbbJ
CCtdD2WwEGn6areKvJoUcWT5aV3DlFBAg/pSArjuQl3SqhAph4TyQdRtTH5gSa/1xJAeYKnZapr+
aKl79Tn7zGwsEum2tL2jcq3gWLRVaQZqoLdXzBMCyowqBxUXvi4xUs4hSYI1e7yZmBVFdUUNjaQS
Lm8cKkFDvqpLsxUFC4xwJ6Qy4nE1CUn/pjIBHTZcUgjemUAWu4MK/6lRuTSYtvnunyL4T54ibZHj
Sg4MSXVenLZ6aUKTkKc2WIl+LlSDlfYK9ufnN5ceWw/6trfEZ3GPxYlYOqBUEGp7E8C+X3gQRDh4
TT/Oi7dknD10fL+SBN8bblMpedADjDZ9FVvTMe4eMcmOLXx6Du1HK9vjbI4/zt1bEbv/IXI2Wygn
m7Zc3UZHm3AyHxCSgT7kYgjGE1mOxdOP9AXT0W+bHhK7mBqeX1/CHi3rkVnTmGgpyqZkxwP5+t7b
hTF5ucaDiGP9kGUXIxqbINtAK/WVd2+rCGy8ESRdldnU7HMxeXLQHA7qDN3ffQy7j6HlQgt6JZ0V
z5SanH76YtLoXpoBJu0S6aQNbPVez6kc/sNw6qQTUwqnG4SmyWvpE63S6jETEKfI9NnSTy1Z9TTz
s8bTUdEQCpcq8FOxWePg5WtZCGnu97zys7fmtF3uXvxDFC4KGmbM3bzCxs3VgMmVABM1UdarMMV2
nDKm8QHuIA01F5qBWuaYMENXgT8FBMxToE4vuUHI63mIRgCM2VgRRoavTN8/PpHRKlQIWvGJS/I8
3a3cdslB9pQMlh2rURM2kJ28C+amTyKR2/9ajkG0vWX+aPrO/LJm5UA0DyD64BRBtwTZifqLP7Ew
v9L1bc5aT42q2rNawHVGmWgGPzbY2ay/2lL/F3lLmyQRDIzFk7LECJE9H8clYNA9PzK5KBbgrbbK
1iOy27Zstg9lRrfGAn7YU9u4lFGqs0ZIlSrEAFdHgI+PFnSjWF15Ci4oVu2y1TwI2zTS/bzSywlh
+rWp7OpOsYquZIma53QIUe4aCzY+kv942PJ/KxNQfhc8MTzll7cFv4qkTdo7TWAskhlXUVKMHq04
h843jE+11iS8V7RTYexmk9qepIfohqN9ntJNgwST0ihP6r7HCwH2fabD+mh8vMou+gQnRot3KEgQ
vdxU1kg1AYPtqJ1J6o9ttA12cM7dK5SZh/Zq+btms74enYktRuaNsEUnzlf82eefvk6/J5bIAJIy
i9R0a0iOFVGe3jSoghykPaw4XMpeEW+KkbWwnyMKrMUDeftgGGpEvQdaFv1ocRwyiBgehC7nCKaT
XFsht8a2bdk/pl5uZWR7VtBX79Bj1p8vNX1fzthjsrao/FfMmo8twTdEWn71KrGF9ssfjkNDX1s+
U99NexTso2/TdoA/ckP6g8/zL2tYvVhjDSUzHo79G6avUpdFh1NxkkoaSIgh2KwtegnBi6BiyFSp
ohyhDlWlJkq4uj3dF8ZqjBwCl9CGgZjbEuYcxXyBoL2p2S0OhK19WNycsJVtOns8Fi8CR4WgG9aJ
jRQt4RvHFk6X7SfkeSTGvCpqXOwCdQWOearwLjd3rvwaWViRXu/wZImFaIRTVNvlTnDuUxn15K4D
AxZCqjnOp9XTGogGUri1rmtrsOJ6l9d452JsvfWJIzUFMTz5N6x5SaM5mTBojV5UwiilX0hSFocF
+6YfbPlImff9GrEB90OMFqk+TG519JiwD/Q2GOFdPOleIfQ3nql9Za6rIy4bL6ooCRS+RBMCGRFO
4I43BOqmcJ1U2Y6DvXI38V2mCA582K+XlJiGHArbWwQMVtSCoHDrwI8s304f0Ev+EtbCc+e5kHls
OVroWr4/lMWfnpz+P/WImP88v/9atUpH3kfkk8F+2gp1KenXpgLIVKXXN4/dDEiOrvr09emjoo7O
MOxj9OFAREMvWOBKdziJ8TxWD9YCkr3HjTNaLn+Vp4iHD6wXlVjokhm/g9NJPOwGlTmHlPehueOZ
kRTWpooHfENEW1H+ucxSfF01SCujpbxxvC0FPoWdatjJvnVEefq7EMneDhUlhzsSAHuSUDl1R7Lw
U/iuRQjk2bSvvxOo0xLBsz4GiRSgkQVsCxmDOzD9dxigwvfJ9f1b9F99Gbiovohxf4sqrmKwVumS
xpXZgqJ55YYpqExjdJmVMaAnxEK6Zi+6bcJaobvTGQvWlg+2+pGH+3TQTM/n5gKYtBMGjrteyKb7
8hvwQNjTfJ0vHZZVXiiDowncMvmSR4EDwf6IPYR3KR3KLCIiEygP+YkndEAksW3RK4gRUEu4eew3
0sM7otZPSwa5+rRSHIrCx7g5iftjhswL0YhLcGbsMbNRF9SXXFPATgWMlhECfEIWcxOb3D02ir2F
IX2M05lOEYXTCOtMXJMl7XDmZTW+KfrVUqRiVJugCQM563hcYqJDBNQxSyy7n0D3y1FnHIk78lEA
FZDdn4dUnJqvnzh2gNkn45O8G4zUYfVEsRDJkvZr2PqQcXbn3c+tjNeThqKGEbtQEnmZ8io43HB8
FqqZmTb2t1/sjCLyu6qdIP3sToev+na6vFEOfthtl9k3YltwF+UQrWXZyO3Kkl0QsEJmajlTu+CW
urGqiNWvj4nmoWjaNPRzsKjFUVYm5alD5Khbq/EYps4bk8EZEyGo6cmqg7Jn1gur2EmrlbPXacfI
weTjOOOWdx5lgRCBIfDXRJmfYFzesfQy54hSQIVX9ko2DKOo1J31EwbyIvrQo8+r81FbdtNewi/L
wUEdBxv+TuzHK3qdMDYyMUvX9x4t9/tW9DdVHgjvE9RSME7dWIg9PRuwb1/aT0metWoYR4AyDNco
nbyCBXCWcyTdI3xOmFIU6zl0doApuqUI87zs2lzjxIk4j53rdNY5bsY+lNz14I2YRU8weM/MnT+P
wEVdqflZ7JSdJILq3wAMzu9jOF4ouCuzCF4UEXaYAkRHUMX9Y46BYbcwwxCL6H+2+3v+Wsa9xGOe
xDVWfxqARQ4aw/dS13RkeHbKg2gc3n7ukMZW2X8zAWaWi5ca5lYw6BxLcTpicAYMtfMUT++oLHpl
q0RxNs/d4RfiHqty7c16kNwwgRicKvN93rKAzaT0lTZQ8hvXw8FGHCGEPefku6hiemA29Yzn9Eb1
st6mANICXMYKckEG0Nj6U0G60mLX5e173juAvPPT3hDY0JRs1w99uGGRBCG5o3QPk4MoG6fMRI7A
vbUF0POrH6w4nH8EnLO/dK3VgUpkzgl7YmcMkLEwOFSNbvV7m8kK5VVq7MVBbWBHWochVzd4ZQvi
FSd5Yrtw4gBqKXTSA7nBT4GRvDEiQl06f1kLeat1+xyDR4SF18ryfVoXkaBsKdlw7Z4osfs5XOz6
iUnZv/ZETklwP7ZsmXDqgQ2Et85f75PZ3czE7lKXMJOcIStSMfTNsCoid+3O2dlAzu39wDkXBp3p
LmWkylciYfk+hiwo1y7uWvZUguYyg6V1FbUWNXJdH+w1iXp5P5ROoYUrA+JE+xVVFQW0bZ7itddh
dLz+fFLaclcToTr0rcrvn7wd2jewcIdo1+ait1YW42ch+dgKY1QhEtUJxwdxJVZVtbLzB56xbcep
bXsRomdbd2+Y5pkGI5Kq9fDJNetUZ6grs9ywU7hx3ORIkyPieR1VJ007BzfjwNpxkFYoZoudib3A
+jdQKWdCOScprmgTmVwezL1XexsQ24u4pf9xB19Kuih1SRLsOZ5PV2etUX4yIIsp1iUbJ6leUhNq
WGPY2vdw4oJCANd6RbXvI/OF+WZrYxZzmotpGrt/sok545fMbu+9nJVIqStRQVILsumd6McVG2ur
dBHg/0Opv4aabSQ8akdh+NB6kVeaFWSjrHdkLvIQWRJm9Gyrf3XzRdscDr/PXdagsj5q1JaoKnEa
F4Zzlq1lNXIyL+w/KLYJPNbHHy09fp8waYkQUWgE6iQQkSA8DjQJO8spivx/H7ZC5zuj+2arpXjY
G+VKrd9Jef4YIPKy362a8u3vpWBCeazvxDMTosnPYVPD4sU6WHV2VjodhNWWDM2npm0cvmx2lQPL
SzLH2vuUNa96K/zG1QKyAtKjsO2OV4BUVXpp7D49uhG5sdU+MStPS8N6gWhhhETJs+fTS8a4odAq
whxVpgxBPvCyuGQltLcnAwskf575P/qMVzIcMbqKg9CWlSgxHLdGhpFX4D3vdec6XHe7JJkAsB8D
wYxNpw9PgSnSf529ZJ5bN0OwiBCevoEYixPjY5AoOz8nYOovtBKloZx1vJcy0n1dKs9HrqjgsmoW
moHW5r6rNHD8ASqW3woKwWFsJlMRMTR0VoDdlybsQokNLe96wa460K034WbzRP8VGD4PgVrISRST
RPmbLSR+YRT+PNtWMVs+t0DIFeSuEVYEYrHoPBYiCmJ2kZAXJbXkLjkwbZGtZcqRAopsRtmY6ZHO
jAERoNKHsUC68tzbo8Iq0UxQYDnwLg7zqQ9qiaEXRsgTCdvH5W44dvLwlyjDtUryX7qXe74q8PvU
eCPbdhEYEoAkkPRqsXnfwJHDH0RbCK0dBspXT4zMW+EGGZd/oc0JaXkcWisOoYIgmMVE8cyJjwem
uPsHlFbdSq5rVU9QwjRehYFavBcVYAw+sS2zNGQHKRYiV1i3FPXmq6Pe6D/3Ylfnxs527FafB0/E
zVT4IcsQfC35sqSn+sTQr80eP2QFy46jTJi9Zh4J0c/0zk2hSQSJnephscRJJMGi0CBKraBmTpTj
U/Ht/heNPbT8CIQ/MM6brbfZ5KI95lB96FUgbrLWv1vSsRirMBXRasPQfLXsUn2TPZuivjEn1QXC
L5wqgtGFFPLrWIEzCT5HtImjbmX4jCkj212xK6ABAyNmBtuEulkug+2Vxic3uTjL90hDlqMz/pJO
MpIblcBPB6PHAIbt+uAzmmM4SnifSySNS66mi+nj2PobnMK/SfGt9ab7cFUXRKcjyFKSd2V6U6tn
8NGjgBgAnWywepaHQxlYkqYeJG643+YAb2Oc1dYAyWJJKWOpJP7paTfdc30RTcbUDYW+NUpf4W4I
dLGUSpjZM3GbqIHlQPX9LKmPHYPC0l/w8yFwBJNRCORoplkLhlQa6M/F9UrCqdJwGq3YEl7DhGiw
l8y19a08udWZ/dWXjQW/cZFqTAqEHv/wNmwULu6tiZkxP5Q/GXBZmEefE4WgakdtgknR3nYJGd2l
ifCdsBatp4aorDqtbqTSzFXgtCRASDYLTHfxVZz5jez/qN5orbDUZnmFreK0+/q/0UzOq1bXxSw/
4jd7TcyIrFnny+U6wVe7uL2oVoSsYj6NTgMXPWtLVpGtmBFszetSZSnOAL9AYF84LeTBX7A1erwL
QdkvXeHrWoq55XFZsrspLIjuzkF3MnrMJXtalGrkwIiOq9ICCpKhRjvnBhYfjspxhR89gd2p1Tkg
VzACUrawjILVb5Bov+xlFMpXT+kLmono4SwkNFy+DG8aS8ACS9piRknJyu2rQHhLUhJPtaai2tVb
6tFCd2SnZ6pSywYK/mGUSZzgKXHB78Im8fzKIOTKUjAx2CghzRjPHOcQlZIIB/1V06ICtmfVyvoh
+eRFPI4kza4bVgVMnvGSi36DuwN5sLwq9WHxemlnnvbilwk1TybyNd6Usz1Q2m0V/vuaT+KaOQsX
pIcxDWaRbmhWj0zhpD3rUTBF72hAD7x1OkMF7hDgRsyntykpCRlAdITl8Crxt+mnixCImTfL0j4E
+9PMF46NS05af1xOBnLujSc7T1KDZjtfqx+Yrzk3/lN/qRlaFVp9d9e+eWjijz56WJwS+AAsvMkQ
VgU8G+u2TWKanfGrbHjUf9c+hu7V9TJIz0afiGzLQ3D1mJmRwZh4nVgDhUuaQoDb4I46UX4Lw4M1
yXl6Mp60MdRtJwy3SC4RweX9UxRCLxeAfGiI5vT/rNA9C1l5YbF+MV6qKE7L+XZAOU5kDZ7IcP5p
RoapjkWe3BuI4076fc5K7gd6wKlHLp9B7r2N/iBc/SRFTolPF/TInxAG+i23bbCy6pe42axJxEta
mO468tcrffJoo1RfOP35UDq6Gqi/tl80UVZB+r2SgBEDCNg9+4SdkZLC+/bZ4PkiqbZ7q4LH0WX6
fvmMPptJsmKM9RjaN1PIQtyOKlIce4emm08wC4ke6059fEHInjuYGlw3GFCkE+iWFDcxeOXCrtVC
WFUQTgHTzVMyR7CJa1Twhjl86UprFTwBf/GBWnktdwKfd7iNIRxT116srsdbWDPD747zK/4EH2aY
QQ0+kSIMaC10q9Qu+xleQJnm66lfyS8jktPn7LbPNYB1noD8030mjWTDSV0QMRoAVo3pUNjMw6UE
4PaXZCGo0xDC2MJsDU/mR2htK9B65aKGqgxnHSwbztfEVuV5rqD02sDVFhsLSPeidzhvidOU+Rb7
0Q/5xj8q3koBmcATAuR1hG/kuQAd6zw4Thxqt4eb3XXJh2A+KkJ9wu5j54gOkSFmerJ6KNiVKtyE
TMdH545iqzmuCM9Biyq3l6+JDL5OKGcnfCmLCKyppT5W67PKszkFisjsI5u89I+OWGa4PX6e4CKQ
PNEXmiuSTMmzAm3C9jg9LGebBJfPX5KqBU9slekwf1t2+zWZCzpXqiYVwJLqFoTya3ZK8Yjngh3C
zCxM/Fsmfi+e2/OOGOZCnGqYrS+pVZjqlX7Hxp0DCd7ZryFIF2L81gN/vCqQBlruMe8OOW+xzpx4
5iZ3yii84bqpjVtOUdQBjSRTzf3rsRhhKh/dliVezXzLoCHdHIPMiLcrWJnOiKR9NAEKUI/5+YqY
l8OlJZQXUN+mBesA0cPcxvC9Dd5turo6yTTq8LTee8d8rgMOIHvAIBR0ZbDhJOzBBTdqsKvMuLIs
9A4Qn+NoJRiN6Yp9m+YSF+YjMP3IDrRBciGZxECa3zjDjH0Rkg58Vw9h5Mo+UFT57IKnGTY2ApX9
mW+jsm6HSVJIAtNGdKjqYxs5xaow6A+WveYJi3DexFaKItDFI2pcEryUxIawm1VHs3klzpPSKozB
nJl1P3lnKfvAO/bUBWsmQwgsrt1brH5Gl6g1zw5xGm3GnG/i7rBl7e8MTSFpa25KCgDKmBvliTH6
RfKSqfRQLeZxV8P3zehIG69BYmgccvnbhj7SGLTGwtQkLjfqazGPYpBq4ringa3MIaHFj0fpXqV5
LsVrNiSqrpUwZMu05v7DdR2NtEpC/59YZt93xQ15V+F5ByJHSRrORe7PzybK2b7p4Hr2Z4MTiGw8
BaxvyLKDS45Fyhz1Tx4LYDrmDluqLe9SG3XgYWn5AxoEfKVDfh09Er9UJ+CnxAI4dpd1DO8Ci+3o
/7JK/Q0hez44NPMIurxW8XefhOwBHOW97OywRTj9YRTIn0by5T0XLd52R+3VxBanZSEOHMSVxoGX
x7LiqJjjLkMhiCrDgP0zdyv56/tuK6Iq+8fb1c2HzXdh246qzkA6f9/hsRv5oHLVZ767c6x5v5U/
D9OC/wCu5mSFYsJuYl23f+N+M2/EaDWF26scuMBIeCcDIsNtXQF3l1bCz3aoJyLNWmZen568ikWI
x1LIQcCGRON/wD6+gCwErm+OzdDrQuUqsIy6bal8MRlFcuPjGYDNedDhIk5AKyzGH5M3VVEbSm/m
B38aCnSjq5s8+zvGu29Ht93JTDl4g8Tf49oRGGOVjzqsrwsFvZ8lZJBXvQHoOlj7nLmflDtmRU6V
WSHJb3jXMjAN5l2gAaIcn2Oq9qzbVUEQls+IBB5q6aLtfqiWRbw8mTgI2A3UxL6uEY0qWXrJckKe
hWXPykybLidUjVbT3HMPIm437Jhg+lzsmExPK4SaqaZDJzXDhKsYTmTZjusUcQG/+A+A6pNGxiyE
psHmuhIw2KVCfDQGUKtEZVArbXabvuzSNOk8T3/L9i2JGpCr/hgLXkYZ+68d9U/J9efiAoFM5wjI
LbM/venVKrBroUrZGvo32k/cknXW+d4G21x1OIWP8V/v/7YWyFzUTnkQLSEeee8jJlubSgFu1lym
dsf5CpzJg6tU8C76EXeeBpCws0B9PbaSRngnRuxoeWSp65cennMh3yVOPAJHaH33DWG0PhbHpnTY
wnJXVF5vHKbhWHSzgJJHRDPvaTKAClaurS+OuV09MuJmIYHBsYtBnjHomFM4vkoxcS7/ZG+ZiK8z
jHVghn9lIWY3PpvJQOAegqLMH5tLUtQne5BXSdGIAcWL5HgmSjkhS4SV042AFJJAJXnqoKLIss/G
v/Ai3RfX5pmBqXEU8J95c0pCImSDkuntnuAqZkQc7tFZ5qJ1edVdspFXBjMv6EoHPoQkFzY0gqLA
+8B+xx2++97FycG0ePa5HKVQiamXDhe30b8fDxERxZYJCe6bJ/G7zEuSxoBPd6X1UGE9VFegh964
axzLKwHRsewVsRMjWourM9qWpZ+mYyzGxbptKZan/YAW3f1LIne4i8MrMHeN5TcUoVxzsxyaNjFu
Emm/tyGRST68k5TkWWHok5kFCdIaAKQdWoXhb9d7SqSyaVpDrRKwo0dS+znzXPMjTtTQqJjDh5eu
q+CdjpdO2Bodjy3FMGVLSV+jfInuKyofOTlSri85XJQvqwAqvtbFXpFCDpVNtpYL6Z0ZgDapZSJp
4c9+1d+17p0IQVTxhDTH/bcxJLI3fzH3Lmu1oxxsLgAfJHBjoZnkPHZxzGL5xhzXCLZsZhgqJr47
XbYGlS0KBcQ6uMDVPFqsuy4e58C/0x0bIKt2TIxPB44XMd9aNdw0JjRM5xBWMU2tPE2BcWY8N0nR
ghq1c7lStyc5bBFELboO+EqdCwJRQBy8FfxctoCTjaP6ioyJfyvyGiw0gOYSJINt4u0bmufWDCAJ
xIam1bXRlEw+dpTu/SQjxuFnB8HrUH1wHmRfCXLLGVDwtPgJOIDGaiQCdc1fG+KH/GVe/5528e8D
3OmcPnL31dlHGBBq2vVClEcY0lFBv8s5r+GwvfmHlCnZm3SZ/pvIlla2lfoaxA1zHjNgnIvl4RXi
K9pFRG6M68rel9ZGZ6JpmqPF8VV+8n8BZe2uEPy5yPf6PKACxpbDnYevLxbcTaxcvhUd4XAvBeLT
Pg+JWtvqavSt2zd5dZnv7fUMTZm2OhQiWalXr4BhkGtkEGaqdJmiUttvzfb51oKU+mjh33cijODH
pNJJQ880v8aPaB4sq9VkCHlF73ItMuto6rSirlSiN0dvDfgQb2gx/vlo9leYCVn4Iqglqvn84iHH
5LnPaGhc1776WAZ65BqRAnE4omp/yyFlAtYSFq3sxazYeMeBHHmmIfhnqJzmJvNowd+N3XruBSJe
BMGQWp/AAXcXuGKkWj0JcCdUMBbWBRa3mSF2bTkmI5gVuappgIatnqpii8yQX40IlCPAiPN9ZaBf
FvYsMu7rwftt461CZmp5n4sy0E+LNl2CeB70WaY61HOPCNbDzFEyBnQ82UXy/rmSdOFj9m8tpEEh
b0KSsBO+NhKrOMgRROc3lo81BxEwvIhLwd4LQ0wQUBmkAgIaF7Op6wxYlVOqMuwWj1e5dLoYPnpV
yrriuI3/qFuSjm51dMU3r9uFLv1GjkwM8rBIMZw4U6QEvBYOPNsfctd8EZ2iLtrVZeRzS9ayVSG9
kJJJgj7kFXRmvdF+snWJvZZCB7sOBmBB/K4jKFwXh5d84Jkfz+4dthjfO268FUvql+o4Q3HQ4zu6
911I/+u4ROAqSvimYsztItZAxpu/OCIz8VDzMCcnDFPIs6H3VZDDcD62wddNTrndjwTp7CO4e0wb
Y0P8cVoJCnxJPJa2ZQ7/gaRalaEaOxCEqcokqqEL7IUOfb9MeyhcLE8O1uJGMWRBfVDFzKa3OhQF
ffNCvO0uDjG5d1yn/7yko7rEe+66ylcwiS2ScBaoAFR29epNCedkG5V/7qVJZPJgNkmUoSgUNs6r
VecNWhA4IZFjf5PZsi80Ivz16/oIUeexWsf5EnPANbJAmxtI5loEm7DNyvH6vo1/z7aPz+PP1PRq
OUGHC5Xq+QiOCShLtKftzaXSJg1I1Q2aEs3BwH1vxX+KP6I9OgicGOYmjKbn7Gp1hsOHH54T9Phq
qBTMMtm8hI6tEXeTpuuOWcziO7tazh5xlykxb5ZhhcsBbbJ3XC3nKmIUWg0i5CRsCmDHsX6X69sb
+x4yOnbjs4LQPNPKirJKmtg0KaPPytxv6GMFRFk0RU82Vcw5qDgtqKHd6DfmXnqr59DKwipXBeK3
dbAe30vRu7v9GhLth1eB0IPhY5HTWtCz1U1OneiwaE1eTXsmGOR0XBWMmPJ5/CHz4H6i9whrB0c5
pMosJsfhH3Mxv5XTxFDf6DhlRhfN4FcWaW8I4qynzfmRC84xrugPuQPDbo97fB5eCX4Vd/PcxFog
5btZSzGb7ChhLQ6FL4lW0oeEj5hIFe05aWen9kIjhPPbWBbpZvP9OfxzZaYGde3d7GfD6LIDF/hv
YIMOJ4QHi/qRUGjrpNzGYsum1H0032NOh1wF9h7f8fRYx0gzLIZk4Vi2oAjyYx7FmD/T5zJZ7Z3d
IGgENIErgkZsVjXQwiuy/xZbh88gvJuyEX7y9lrGGvimpD+CrqmPH7f5x9/G/uMJzbKgYSiRG09F
IR5izYJzQpJU+zuijvVnPe3yF8IH3PSkBeJW1a5YQ/36E0Yd8Nz1P2ncJ7UlgMaJ94NZsYDEXrR+
KcqqoFEwDQKPdZEZr3mQT7fSYA8Cz7xieDGPsPtFY03/3haBwvkgPXzHRZvWOipUczZVueX78Tto
OztsGTbW9je8sw4zTiuUZcDNk7XLwCUojlRdYxFCEGok1eyfuqKz19Hbtst8o09KOO8rLJkvekoD
5oe5haAfY+Z8gJJ3orSQ/53z6yBEVQ8MBEk9oLF1WnTGQIBhfFfSojJvFomo/HyXdO/mj1hGmHuv
7D/nsfbKwBOVe8A3eFfJhYOxNBnIKG+rElcXZmtE1iPOEaec9SoOsJbgWKovv4WbX0AWF3Kz+AEq
KNHaQkorDQylaMXpzyxETa/SePAesumzYHGE983wddpjhdnf2sUGZ8+bUbfdG00hKJ/6sFfTMaOY
x2mFN38RAMfSjOjbOub6FHb8VhgoRgdsMRFmLDy+7dE0Bf/gDp+z+9ppuzHg7ALMzIvvh9YxxDyQ
jQ0vC7VO89GjXPH569ImcXbnhqWXwyCqP8QI0CsKrYm0qiR9NSwGRLmqpXNejy9uAdelNS8FAkAM
3oZa+2iGPcdqXlpIcd96RFBiPc+kJnmwP8XFObgKvC5WF1MM+ozw1zSnynlR/OQOma7AYsIMVqps
IXT1k0STF8v416WzKiU9QVZg55J4mNGAsojp0f5nL63UPKgVRsz49YmD9dfDgPvEiM46Z/OvEYy+
TD/Yf4zjeSxWhWPN2K9i8clG+7Hg7RALVrFXqvD7nbNQdjbjEK7xZfDnudnoe5w6JFl+6/YTMpHx
0PlvZBjTcUV8fo2Fdd5Ry/vd2AM+MUu0wwA3/bWbhOE+tppACFHpomrapK74s9JZcY/F8DJexBxn
U4H47eaUQVahOxU6QPki/VyRaqr+52NDjZ24BZIIKG0+huXKV6BjQaAYGWoFGXm9VchN+Fu1uuAb
DKetxi9QHAi25xSbqtQDDaI8QfI0iGFJhD+Xb3mGjTqg8YTq2+0sZV7LPVPV+4MMQ4Zob5phkEHX
BgmQEDdiU+PpC1rZ34UGrAPoPI8aSosYU6Cynggr8nvyfd8/lrsnX1Ik6a/TZxfuYZTPsXLZW3o9
lOGD00zVexgyjKoPny7MFEXhC+zlJDVYXnZ1XzMQvZLc/iFlM1u2evDdgJtg8x08E/xs+B8VyuH3
uSWf9eyzDfvSvGLgHaxA4vUYsWZ6yLqS1YUHVXsyDvdUlafO6M0RnKhS1oRMNQIG8p8wOJ+tQVzo
qbLGoqRNZ+okamNwSuVqcvwD2HTzonMVrIzYqlKSglPEp5/vR7uIgu0R+VHZ05nTqtVYGL2mFOTA
RgdwLgFetdteBnd9YyTZpFCt2qKezO1TPfBiyi11sZebm47OxU+ag6p79ffBlb0B/e4NdBajo+gZ
mSprEx8GkZJOPaULtdi1W8dwppzkW+VXFNZv58WSecwMqqGAFWzG92EU9COwmkKc9tyG7mD0mlv0
sAGTjPGhrWkzp7zjmGLxMVHGAb8DlIU3KwFxDGOi9Pgd148g/gH9PwopoM3vjDV12jX3Ije0Blmv
Iug937aVNlKbZ6wvb+DyBFdIbVu5wrisSGKtFnJQ8rdMo3hmNi1OhxaMbcsZIOZc3ZkEN3xyuKSC
fVCoOs6AWgg5r14j8VWCVfci+CrszGv+PRLYRyvimcHF9vsTBaVu2HHj/8pPLEvxes8fRPG3lZJC
nmvBlTbSJS4amCXCRJue9QIsQehisvEsltR+F7x8tJFB86dl1NHZEA0/HnqvpTbJOBS7xzEcAG9B
pboHNBHVyALkOf+xgdo8QX5/+W9G1rkaCanpgZWc4G4FxTsL2tyxE5nhOTXlSh7FUI/6mOoVsxKw
zWG7ipX+D9rvUUAHN3CKxBB/r8WzE8r4aeKRBScxHewR0DLWSgciDMnHkOyR9lY1tQQNkL3v2VsE
jPFYFEEgUB/POka/UNDsx7gmVYccaFAL/R/2PdosPuWR7em8TK2lkl7N4xZRPJ0AsamIjAl6dKg/
weYTob8h07kouoBsNZJ2bPcIAWShQcg/lb9jfo/RB5jB4bvhHxcIC2RCWgRTlmHgdSXUIVcXdUTi
8ZVQ9XIgq04YDqVrini6DpPzRo433pI9TPd5zvmXx3EbZKOrQ02Jl2RCGqWBra/4cbcs3nbVS9bU
JNcWMqiL5yhsRKGTQlmJCyw+GD2zY6xbxUXUQVVM6OzmvcdIxAxOKVL5E2UMkcmk52i0fbOArkzB
KVSCjJ+RM0AZHRzzXzF30Joz9oRpgj5zeOc/2VakXHoXyb00kjgJcke3yuc3Y5v/A3v+yqjoKV+B
xlgk4kO5vaC1l4eT9sJnVN4GtxJEeuDHtnn+ku24JqLC0Occ/3UrkEfJwmfDgLmcfK1ULQ8gKFnI
MzjqhuFJbQcr/PBJ3v+kjrSTi/nX+6tq2mZDf4TWidhpqHG4tAj6Of6uuAbLIGNz6Ai6EdmQKqV5
+wHZw8yqZS9kuSqcXMFnlEgf6GJlUxK/lJ8UgbRhdwXJIK2NhjC0nsFKPDceDjMgxW+d2beq2Cpf
UlAxyje2ZbVs2etmpJ/wjubipdZ9pJy6dS6J2DabCgtjEPXJurvJAO8Bria7BFmv6A4j39+4OtAt
NhPO7/EAhYDo61hEkLo4AmcZr5lZ+eE398OTG1QkR0g2YIIbzv9nh+RCcgpMxeVhnL40O54RZuRK
Cn9Ilwx463uVM9ZLMJl5BmyePjnCNOiY7ABDVcUDukv8wC1WOIc3BF58VCjK/dzLAY+sMiTBrzyy
c/UqTJZNrNWfaD72qR3uOs5mP4+M2qZ7CjcmX3JdBQs7HkeoMkwkfR4G8hHYUdBEk+D4rloy7adc
UTK3Qp2f0d3B+s+tavylh0Usajw4DbS+zWDJqiS/k8IN3RmLeEKgFHyKqnKUHAovsfMwmR0HGzme
JfFIF/KthnYS8yonJfGxs1tpCU6gIU73OhPd93zWRGrFi9fRzXaWZ3VEoGf+SGvYphTqdLZNOVFM
+VYLeCpidZcajPXpmRNG/aHT8u6IuDA+CzESS9rwb/OvrohlnUfXmyaX32nn63MGx3pG49qVdwsY
Kloqq+0axb7RTRBR3E4Pb4+IsVEH17WK7OqPZuP9x2VHN7BfoBZraODGKXt6GxQXttWgkv35eTUX
LhsNFl8X2KYtJTolhODUUZYq7gbTG/joBcphm5K5KK+qgEAUxJh4HX4d9MgEvkvWQoxQOG0WFwoy
6IM4MV3MEGjBbNybfPQbQ5I9limwQEE3H6nXxBMfqpaKBYIKFNoTYiiIUa2vW/hef7omXZLk0+WO
3YjDECnWE3NzGh/mwafcoIDd9p1ttn0fimVlmpaSUnH7NFo0KzbBS0NbRSTYgpn4UPi11Z4iqkyK
nOnykzzap3XVXdfRCek9jc1elXcghCWZT7L/XVSPRrjSjCIOk9iVVwOmbXcPQNpRPd8VOfSpFXfi
8i41yJNCpO58SY/hdMc7mbnLsaym9YW4hicH4CVscU41JmMN0M/9zKT7WA5jQFGXEy9vqDAtn2/b
yr5e0KsYMZFiT3GS4oniM0MAXteb4raY+ID2PXHccFMHgZV4flD45f1N/sXPqi2+2tyyQs7UBLqI
BXhFm6NrrN0jHDl3wXbaKGNP9P2bkCNsfgtM1/H2kxQ+4agqoQUTdvppF7JF/2klrRzSjUSLB2FX
JbICpq1Wgt8oYUzPgFCjnN0160F8vwq/Bd8iTy06QdsEOycqDMteozdgVChvxI8rBO7V9kuMvKXP
FVgT061if8XllpK+EG1vyWklf/LY/mlU+jM7JSh4VA916AN5Ty9VimHExg1ZnT0sHw0I8wgr2W9Z
ZCMNv/zdIwMQqndxq8mk+4E9kqcRpeQ5T61o+L1ORFRYdwhP+ziFwIu+vPnony2s+SQ/6qk4re4u
tlLgewYOdKrLBVOx7vctKhAfzykNzhztqlMM7bnC3320Yxhb0igfo5RNcIpGPEjdBUr9QFU4fPXp
yYs5OlpoY7lwvKWTj+klqSTTtH+aJCcdjppxAMuc7a56Y963ylPfY6uAsR4jfHbTWWnQQllXVvtB
5VDLPpLaJ9EY0SR7whTcEJohEJnvFuR/Lr+tJeG8k4BOFtuYN4MLS9l4LiEojvUlWNP/gSbRqSjn
CezHoZBPS6tKQmCAB3Fviv/lKnUJbX48hYMfdqNwkdyyy25uX8s227rhGae0VJOPAMMLZfivmjWa
koxxDOZffRTszrmlb4QrLvOndVsKWgvaEYgUkajUdlJf0/y+EgCns5wCxuNP20n0dXXvYnCT5wO4
pk4erj7X7fYyKMaV9MvBbgzjkm1ffNePv0cEciSUCeL+4P5Gv6NPiJjXVbGiOD+XbtH1X3ggMoFB
VCd36R/1JHRChLuF5k95L6jORIytJw+2WyhK0hRbrxJf8pbHis98DBreBQ8lPa3zzST0K7zb1uQx
bGD8WFezCWSsjXZAg4UtwVr8PC0M+/UIZ+seDTJLsPqF1XBnpJxPRGkaJOZRt+XRlnsdDpUDm8YF
cSUdcVNCxVbWzEnnLStJkqF/jSPIQS1qICyVmOrAv6J3M9+pBAMW9LHnjT/jxHJtGr3yyLaACjre
zodd0ARx/LoZDpNKx7gclyf5GRFHGCppcOiPGnrxKCxAcCpscmJAlvR5AyAIpdUIV/TbcB8FcGer
CI+w73o9t3cPCYA8qLOP7e4mBcJ7UQG3l/Ws01rgmpxvaB/GeQLaGMhlIKyw4TIfz5ttcVdMpiTd
xcCfegSPSyXP1YqPhlvoV42d+VraA19MDur9A9XtGJwiHoN9n7TzSetjh5+l4YyHC41v/zmLOdib
U1T26avXMbTg20U0GqB2YohkYVUkRdh6GZ/1r5rjyQx19a6A3qpfgUb8YUIJVTHSx0b6kRp0WUye
DFJhrNaXuVObBqwl9zozbFm8sxgA/LMyi4E0k1VpZELKvJxgTwPF7ThCabvtv6CJs4qLFDPbP87F
3vHLjxCMDJfs8W0FrqikRtDfNhVp7xYo7qcU4V8NcFx58D0U+84f/qtTR9TWOdLU7jK2r8fppRL6
2rMvY2qrnaaZUK+olTkBxtV7iS9/yDN5wpiGyDVVz0Q5BqNJ+imDiv4RdOWiijHvW2qwrK4HCJKu
jHptsEFitcoAvnk72SzO2SIGrq6PlPJACjmOaREJ9u+YF3wYoTfC4FbaNAtR5x2WGKOwabO1bzoG
rKucOuqmzGIoYOnjyqx15yV95f/DTuLt4UX8A0/rohScgURQlN9ssz3Zvcb2ODnMVvsDjfCL+PcJ
aN/dsZGYR0i5fFIOgvENVVw1+cgX4VWPcYRgf4tWmM0LbAnCExgn72u43ROzd9ya9UWaeAvQWtFC
a99r82MMPixJKGBBaS3RxzdVd4IIlSq1/fjTuGLrYBAI8pPIpiF6RoHiD8R4qxuDI+zBlfU7KWQO
X0836eH1HdQtUk4Qzcoour18wO4y588XLbujfk/Uxp6nxbLgA93Dvbq/L9yuPPq26RmKkSFTb49l
Bob3vj/ZZHGBpUjNAN3Dx13rLqeu34upy49JcF6XLS4OkiUEck802V1t5/6GTtfpULxOJHUrw7Nv
H8pJxsgvp4fOdeNfr5/uFevgnEGF6duH/HmNWn1Wz3jGoXIHJh9blEI7iWHpm7GYd68zhxKxLMPD
uLeOvncWrN57NvTgsaQE7e25ZuisXRty1Z4ZU2ke1gnc6n1+qnJfaa/d774beDJp5MkZWSYBjtkM
sSIoTPrWUhs16jqGbkwsKo0fpO8nqLtGoHw90TptcnkHIgjgqYwfk3BdJk+s9y9y3rodio/vFu1Z
ZFk/wTdaGCJnzr38cq4tRcMq4np0OQT2gV9reZNm0gk+yOyyRBPNS6TsIFLCGHQpYc79CPnSVCOS
UCw3yhdc1NfOV+M56Q+VB6o5ouPWzDIv3HLXtdcDXobV5BTTTkQcgPDJ0uTEz4c84NeF+3iOXys9
Blqk1XhjHlBzNKpAl21zP8Gm3J2srTw6azRY+DyiAdLDwC8FawPUYsOHpjixdS2ZuitbA8Xyt6q1
kAIq3hxvfCCD8Pynv1vUxP5EQOB2SwwgwLG8L6QWAe80cAtReKUKYxqHNQIV6VdJnhd77nC6uuky
Yv0MP1ouH+V/LXW6d6DTo5Yv+Z1j4aKyTK/wvbFPSbygUAX6Hb3Fb1BM0dyV7F6tWipE9whIw2iT
zTisEVIH0ZaUAFuLKztRcaSUpVTLdQJwlNh5sGx46jviWHrXW6wrr0t7LqGP7vHW9AbuVeQ64ZOX
wMjCYSyuTPI25JL/XPKYtfj9hJ8UiIyAk5stXg/JMLA6G0xE5mOtye5Au7KxQXHLizZvIA4ylxhD
2rhMVmqcSpeAuDN9kWnhNwh4eH71l2+Kr01mBhA4hF5X9V+dbYZC7VGjTliHdfl6MSTXVPObkW0D
bIZcPv8icmmGdn8mJ06nWXI3S8UBLXmOCF6qjWw68X3N7sICCwiwomgU1UYbi57ORnwE2V2kZSFF
WbWuzY0gJhbaFgvom9AasAzgqRuGjn+nVWPeN+Fk0j07iOXsQK7RTzCLTNxF4GzLCwpjuj0vEA18
Vjokkw4sm6iofMF+YbUjxYYr+oTXyEU1snw6gMH0fpTnM56uzld3mBxj9EYqIbQBI+G/3GqYavF5
MaSpVHzmUy8zBr0+R5fIV8LgHyS3xQIZljfyBZ7HSz2amORhew9IrIU2BBCpYd1PlKzVY9GQWub0
4ytGzuulXTu7Th+eZEIswKIrYte2VmpxtB5wqILspzBngZueaNyFg78h1QEjLgMCdq2V6VCoTPLx
ihQPS3SlGPZybXkLhNzpqhdGI1JLhNhc8xCN5vL0JQet7AWETdyy4JdUi9cL+sGzeQthcY878yiC
YmCvD8U8B2CobDeG/4YEAh0L/qo3hvOWBBwyXAmNkYJqO8iy8dWMSxA6svpOIQ7I9sY22OL6EZWu
cjSU1lS9EABD/se+Rsq7FtRSgpm0NKCDF9baBW1XdVKBSD2CoIcwmVqpiHI6m4rsoLhV1ka0cqNO
or3nH4ZvA9XDK7UKKLyoyO551slEq939R/MQcWyT0Uc5Mgt+QzUgK80IYPLPfd5yOiEeFB8zUTgY
Xc15/ISKwXKaSZOlps6d8d+fP3GE7cdXC7rShqLkTmQdTVlocyyM1ypHnTxpLOXAnfWPhC1DKmD+
1LaRB1vUzO6zZV8bM/gs1pE9CoA4OIH6GkO1jncBz/kDsmATS5qDFIflmHbiZdmzAmVd7UDWQQnu
exm54TKOBF76jri14g80ytDk0ZpjwiMU5u/+UoPSpB/MEaHw8R6VyPV8aZ2qgdqI0R21Yd3m456s
KRLbuVcfD01F8T6GqbyTy5pDoX+bhovn1F4RAFUMDztIpo8mGhn3L0QG9Z30a0j73yp6KbJogexu
oZ8L4saZPQnvk9dHtVr4CrqUyN/52wxRHDFDzL8UhllINJg/CR6RV80J2LOxx+kc2JDktFiq/qFH
CgFHIOtBdxTukQnJ5XEaOGve/eqX5QZrJL02eOzdeVs9miNdYRr5WFixSActxMP6Ft+Jrx7IhygZ
aMDynDwhD2tUuV8UmoVTj+fhuzk7zEMEaBDobtHX/zrJLQadS1PK5twBStSTNJGAc1cOXXwKktB6
/nhoDBlWSGrp4z4TIFziZVZCz163vmaI+7opIfL7Y/e3dGIBZT/bMuq5RCHzM1TPtk4VeWAe7DEv
NCWuDLIRbuPenC4NWLfmySJOAAh59zeVabLs1ZG/p8k4X0IrIiKQtx2K7Y9D0EFdLImcCGRJ5VrI
7p8Spi+fySOr0tU0Phqg5djPAnkZD10szCSPzJpL8IuC092zqy83MCChpLxKc/lTXUoEaI388aNX
AdWmCkjNnf3UAV4rBTA/V1f5WDagk3ScX6JN6333JHIdKVJGIpjqZYMi9xKKJoBnCHxD0PeqAp4x
hR7Rx20zK/IE5FS5f47dDKc9xTFu5T+lANXwi77sXJ5jbSxAYgJ/u3kxkjagcooF7PhXc3cRYWRv
b6c3FJ2q6gMaM+C8Lj34ljGyW8cbb0gK2PFz3g6DL86ULIFIuOShEwVv5x56qog3iPfazyAhitSO
WX7sxuy9DEiR/0UHTLMNwDRSFhV0pZJ6ItyIw0i0jEfFyKBYVO8cOICmUOnLtqYODT7guGHsp+69
1RvenY6GGXMSEAKo3CBn3Y7+kx4IQMVMG4oAv9cAhHPPAx8t8CivFsSDya8eva1FSwVcfcaiFPMT
mw48xcOBdNP/kFfVEE50NHvjtbssuy1SxYfjmob8aeXZJ6Us31I6ymqHxfYlTj7VIJoC9/S9dwNB
RK03hUabJWYox5KZv3aQI5NjL0SXoqE+4+Io9HezAURox1kwnutafgrnutnSEJpRPWwm3b9o+D0B
j7jLgjXwVCHPj9TFMreG4kjRdwzxIU/Wl9zMm1Vo8Tyhqsycymw8wM8w5hvcpfcYORoCQOO71POE
6K4YI8WUwZfui/gM0bnAb+IZGLlYmgjoG64wUDN4ajdQi7CJVXzEODeI0mPYXWvbM2nWxW71La3S
TbVY3acKZPtLZE1MvOJHGGg+fjCiVzsqxBjJPs9CFX32vK1dcfq/4hDzc62gV/sC7IcuH7DT0Din
QgUYOzwO5GrL5ckxRTqpumKVKL00BX9dPsRMf0Of314fAO9Ird8iUpGcXOEQUU8O46oG5/HYkY0F
gkTd/eWurHfyVqkgkxFvkUdwrlprU2LxRAzORCaXG13SV6+zUU1ST9qF/Rw7KN/7XaEGXntykAri
Xs3Gn0hPjjzKfFnE+aP06aWxIn/kfzpuDShvyjmR8EqzBfrbzp5GCyfXffXpGlMiV06Xcv6qJrkA
ZscpLJkJVIduBmhsGM0iJZpc5NNDAr0rIK+1ODTl0HYFyfa0/9F7+mMtexwD3oAAJaMzdrPZ5F9G
9A0vkZ5S5f7VgBOus5UENKBJb+uORAU7SdavDUUhcVmVk/575W6xg0GVc/C6qInD//Rgv1JPgC9Y
A51m4HTcgivsn5IgVc7mFU4pEaszuuixDsxwW2X39ieDZuB79ByjNiFBOHBzF7Q6F2hQxy2WcI4S
g/1K34GYMAZQyvWvzPlyeS90XbmFQ5cIAk2Q2+UOp1adWmqtWBu0+UtO/XudLsMuogHiCtkZ6SnI
STnUNLClcJRMhvxMm++DAJrB+1uvhVQunaVp93wwOTr285EzIykqdEVrHEuBRMPj6BPPZlNEnM22
iQZKfMtpHxdzNb51wkYhX214DVr1GvhbHamhHtiV6/dsiU77G3JGYOe+Hunir8pnPeVyHIC5pxkO
LVmYmmGmIQCzSkeegZWqZRBKTGNubvBbg6SkYgApCxH6o8t7aA4GB39SfAC+SxuMYPEcifpvXo4p
A3p+KJlAlxwpBaLjiJ3EHylYibMDU68xpBtsznBHmz19kmDHKll6f2L6uQrPPtvYu69ukhTMSADW
DOGsgTYtvZv5iRez+/gLWFf11lIdkslwwAuU7T94VsW/sVQ/ZrevJGNAaP3efiSfzxSzWWYYK4B9
zl9KMLX1EWmPlWdnbEs0uZ8rhd0aODNVBEMxpQUxVuRgh96wn59kqT7t7ojO5SRAX5vgMuUQgNq/
e0cOGlPKTWv+w/QpJt73KBog99Uv8heRXbI19QWmCvnvbZK9Xr7yRtbhig3XAjuSMJWd6Mf4JySD
xGZf0TRa+VvCPCqwOLzcFwtflUECADGYS0XI0m5y4lWcxnQ99fe57V2lzFrZZQ2ikn0MorwOO5II
IRpfCQPxBkB8x4qkqvVWjO/HvABbvW0ul0XO5TiZgcKFJIZQ6TuPrg2Ageg3Ehix4nLWI7alySKW
2mEkarfhNtVZHCQ8wh/BY7TegwtBVr29c0ivVKv5btnlq7pZzSAmvkZvdpzfkkcfuECWIf+P1jlJ
YH94/hsasAGR83TiAuEWqBWs3SR/6ueeVTk5pB7WqMaylYbp+kImXjybuT4KPNW5l8GV0q86fvlP
OLWcH+2axWUGEOXjC3kJza08Vxnnk7k5czUtsXRGuRFh08nszbc4jWPwoFAQXLd421JilGnA2zXJ
8uhNsXp26la4tqkYhIzS1rnXm3VbADFNSg2axixPPHyJ+y1bHsdRRUFbT+wyY5EzG7u2i6C1/YAz
sS0BqivjQ/UdvUEbJl+BoeA/LYBYweXf0qjHeUmQj92TjnMOnVeDxpqwZWQInPhjPOg7Ph3pOYbB
W6LzOf8dXGm1Bu3BE+SOOTYKaN3guTOJWZ5d4QucPxkH6wkMUN5t1XlsB0/3431Htrgfxy8OqgHD
uVs7TQSB8nOtxwj49Xw8jdFQBRkMJWnyLXiGiEYljeiZ2PQNa+4jDnVO4karxzQhjXmdE/pe3cRh
1HybF6LTPx3PoRyDxkn/ARMC8IrFJMctD/WrraKGVeA/IlmeSxMoWC7N/opXHcn1TRcjTtnyeDMb
WncphCpaugy5MBA9prer7sVmuRq/b7mhG2pEXXWvSKtXQhEijr5ObiuErYeA8LmEE4ImWQpiNJxM
CBL2cgXU1SENMfUMe1+kitjfoWHFbO9h3yaOq9JPVQhDPPScdgDSSk+M+By+jyWFbdN4E3GPGsH1
Vio1kHq5UEXb58n4lRJXRcGkZ59+DkmduUTN0IZWirfr6CwHKF1eY/548WSsW4qAynQrK5LCGoCM
wuoYTDcDOmX0qaegj1+hmlGpNDj/i+cCePmAB14Ds//RzzTdcdU98eM3lA0MbW1OSi3Kep5ZJvo+
qEWwO7cUdJL3Ahk2KnmBTOYWppU5kZkQ4GIxdAv+Tp8I6E0hSAoQXykgfaQAhf6GOq5AupaBHaiU
+nX79YPjNZXX/R1b0bPZDcsOwAO75ovFc0wfEKnxCFd+7midK1J0/pCoPMpLbW+3fR+RU5JcMcP+
3PqgdAHGp8JM1wvm9yqNocHYDhhvKeWm6nfePPNEe4o703M/Cd+Oh89qBw2VHDYVZlIuzVR8jmUy
W0Emo6fZXet5HoMl6tmTUTjrAOmRMoKXJAsaxFrYnwW7BuQXI/Fb+sDoB3y0KCSYYR7V9Ow5pFKR
ZJax4ERBtAf4I4CNTn/8mpZpHTw+eK2VId94V8J1oN9Ivi3AefWLDwKj4RjqZPaKQeOSUeA4MWyp
FrFU10U0PPjUTBsT4F+SHpaOY9Y74gSx4stZS+RS2EW6GMjSPnXOupY6muwQS9UlwAJbGQsQUOWu
a9Vi5aqwOG7ET6BrIQ0pDx8mdllsE0eUHoBJJwgozz/2GEWLLmWwPucDUnZcAJyVV1rYahdbssBf
tXMlQYn2avZhijYTeztg8ceAiiXRvCEwGRN2pJIatgCyTPRxThneEEDCHMjaMTMH7HjE8agoMok2
75rA/qqk0tWWRLntrFCJMvjvyc2HpcE7kI96LTZw+XuuLvhAd3slNqbgfbWIlzphbTM1j7YvrlQ4
BaGyB5xcQp1tGP8p+/l6OLQzvFliuV+9d0VItgTnRk373t5xJYbbPPABXu5/Ad54FzVwIpV6ByvQ
5wQqeCAFh5oPoKOmzxPUKxFeSfx5fjXfOPOsbEVUCRZY/jpUmtjIO7L+6vSMaHXqp4hMgg4k1cOt
BxCOKrsxzyhjM1FJwXPp0QVPeIrGqGVoZQK+VrQn6RpR5k16jArNQ6JUEaHl79lia6dfKmiOtKRU
dLmP2p7wsUjXu4c3M945MJx3hp2BZPaT1VLSm9XzfTP1+hKZJm9lCk3ZTkkuMJF3XDnK3GAPNUvy
3DlJvAk2p/nuu+VQSPx5jAXbkwR9Rw4GNmtrx6q3CLdY1b/6Qy3o4A3uE+01YUJzwzzSeL/jVYmE
yYJ6KWe3otmUisrPyVCf2AXB19nzwoBic/z/uErfpC91r2YMvzNkXM3EintTX9BcA8k6gnX7dnh2
1vki+KpWbzJlS9EoR4zfOf1vI6VGBdTwLpy+RpgClBWwFywQ7emAskVaZ2ER6e6leLOMLhQTIe3r
kvlyeo0FcTpMhM3S0wclrwt4DN8hivkh6+ceZRIWn7rhqMzH5xlN6OoYeVHzpuuBEZFW7/bFY9kT
N4hLOSbGZvBPE2gqzw2eWLxVlSTWwXLdkD+M13XCQfxyO+a70jeCvpcsuZkaq20cGK56Ilxi3w9i
nZXZIBHjlNAwPPJwc1ZttGrUTGCXuLusjPFEKL5ea1lXrulXLyx2lmSOXvtjnalo6h31N1Rthc/h
9YK9MWGrHgK2p80CiAdLmyZ+o7Zn2wQIiacPQl4GOVSBl12FDZxnqgvDfBy/PY0V8CLhA4wU4ix6
xWq7//7sorPf4u7tMAKZAt6vMO3f2ISQBku7bJDY1QvWhi+WHJF5DSNZ6IrYygmi3ODTKbCATSjo
vbARBYuM+xus8K0i6VYms/qQWVLQaP7s4QCTsi+vOp4bhAiFwthx1mXst8B5krCswQvWbEAbd0uD
gTRuyqP0uV/JPO1dZLqtEKofOin/jizbpaDNiPjt251DsbgQmwCTik3iML0FvM87KecSk3SSJXdy
eF0gmrZC1Brwwg1wr1yesxcgtXN4MBBc/IHn9xnYXnZRJwTjXTVoWkXq88SKvD+XfIFj/eGd7u5l
BT72V6opysTgG4RqsgIjr3D1FsdwCQ5i15IgtL2JMEpWMcjaxVNH/lQQqRn3WHRVZIQTdbDzId4b
QQzaJkXxCAH/0TDZ00kTbOg1aSTKrXvWE8GYOmVm02vRyvYY+fXFwS0MYfIkDeuKsQilC8B0aJiY
jwdscqipmAVKERKD5vtixp9xhC6brvsATYPTUz2nMVUONFpxg/zEQf/WZkVwJUZp1EHVlvzyGuXi
Sw5+QnwsR5xCDOe/c3I3+r13jLYhJabUJNR51FAlCqFX0AZCflLuhubNgyNhDUonju1dLiacuW+C
EaCAIkI/ADrZJORbWXXXCnprqeJdlxfHgKKKZGJ8pFPfkKWudIgZbdyi30TErn3WERxPzWiBxx9d
byBGBUrwcdsgF7UMqRSJ4Wbd5YyTVFt0F1G4LbI8OLHijUbfKKwwpgOHuEo6hm3Sa/Qr/1727Epu
qtHd/CW6CNpEDLOZq/9PYYYipFPlAATGK9HeV6e2JdNU2OVZQdgJyQSL/JiaJIGNjEDeE041Xqwu
LkW+9JvIbtpfjxukk+heGMIcQHBE5ayvsKmmjC+raO0HrjNhuPLD5gK8PipJuBPazAXehexKFwmD
la7CQdxCz/17P7BtZ0Bw+c94ZA5on495qMb5SedvAzfak5f2kcGQ7FaIxBYRDGwz3s2KK8XpF3m3
LE8IX+f8BLz0XuTYDxnACMXWvQKRbKF8/RnoIO4MrC9ofFwE6VW6igqecw7F1G6OZsEBITlLF/KD
0gZcu8vb0iL3ulJFaBa7qXePmodS7L+o4S10RHcG94NUWP9NHXA9Xv+pSMNduBik71eIZmjrvlM5
/7LSQvc5tmBjqPPAWTnHDhTw3AX1g4dlx4g3oKw8y3w1BQvP7uoGlsNiakI4XONP6c7FnCTWgj1S
MVczlQpOgCj1/7bwmBLEr4Ur1WrVrRQsSB52x+JWk+ncqJSBPswmuU8tGyKgJySrOcNVI3wZNS7H
ArccOKsPgJsQNW/H3YhMtXXyB+2ev90410cdX6CDip1gIywHkrpDR6UgxfFPStGoSk6RmEx/IaNm
nkFrtkcA0pgWthq8t0gwOAkOKvRfjjhg651o1J2nTquqP7JO9tn8H6AjQ54NOCn10G1R2XoHjdH4
2wx/16UGXcGIn8hsh9qRt6/CyTv9QlxdSdekHHeIe/vY30y8b/uGH3u+l6sBnsCup59I+CkP6Obi
vtcko2OYVsnu6QB8z69Fdm/hBLuYeFYh6XNd1w7jWb2hF0A7XB1h8kM952cfzxABJnpyAINKH6r6
2amY/TepsQZDKhadz4nmj1hQxxI4o7NxNxookOkM9mZ9ri0XnDelN5Exx2Uhu2qfZ4yuTF2Jx7kB
+1JI0+9dABJ3Dkkh3asomM9Kzu7tBeyizrCk8Gl98AjikRf7d7R1tsgQecApEcSym9Dvyivn59Po
8i5hYHct9eAWHwXPkp7/w38jMeMtTA4/vFFwZL8iemUPwVDF2hdvMCCswc2z2R+JkXc2kkT4J3R5
ibLz8p0VRgPVUVm7HgvgRfD6XBRnwbOQ2rZ8cUcD5oTSMHH5EQzvee7NDINiyZ++iRkWJVB2Vjl1
UffzSNpJ/Xz+OdmFfXHMeNMGhOAdyxe5C0gczugw9e6P9mwdD5WaKuKEzlTaqOCRtGi3dLXnSZ+R
ZgEqGCu9rYKeJ3RDfrcrHmlv5RI6pSh2pU8gyM9HjpfjnxbwTealkHiOk1k1b+6L+vDU3JQ0qam2
jDXsCbHMm9ru92S4ebTvZFWCvoon64vvKqgSvIzdSXX7sp7FzUoWTL3GtXlskO/bfvSthWEOBcZz
C7HPj7mZhU7SYWi4l+NldJNTVXVjUSijlTRghjJSPWATvWg9kRUETv63+ZhIV/okmGEYjpjPLUuw
+UFvHlwx9zHorTCao30imtD+5tL8COHEbLkgbzLplb7AKLjf2/s4PIvXY0eQiufFrGJBokoRjNrB
n490VXGK0nhoBJR+b6hmB784S6gIKZP2AyzbxiH2lI8bFjA9wjdQUH0tYX5E4HY2QYhoeFmZThng
WkaO+WcmbHeucPfgzfB1BHZZ89m3VFQJScAVKghGFKonOgUJJjFaG0SRdanjXcS2PQ2OukjuB0uY
nh/qLSUE97Qk7oKISeaa8S3MX9lW6yTmsRzH2b6IB6rTciENzlLSpT4cmC52rM0LyQxvxP29YsgH
uLr9m6NzlzcLvyKg/jhAb8ddPYbnAymJWRQ/nGhk6nkB/cjQmvXLK8ZDXus4RwMt/FaGDyjCZNx/
Co4LfRGAUF4V23qSQP4rM4n6+fR2p7vkaDgWuj+dmAT9ixnhUI9vrUP6+oqZtoI75zuZr5IvEiAl
5DQOQO2dfLvn1msvztYGuKGW3UzCx3wo7z5KCbI8FIstnUadOiXM+uLwVaBl8zOvVq/RfVSFbxq4
qYgEF5i9/IBk83qRYV7rESTGllt65h6H5/w+1WoWvLrjS+vkg4hbm8sv44kuBgtl3VbXXbjD28ta
O0exYcQ69+u0xScyE68PHn2Ij6uMjN2jjvkDi2trpZBRdmqfVagheVARxRm4UuW83brKxnMMPtfa
BSfYk7FGH+6LEW8C4sWhsSkIQjCUoDpSHl5bBrBYO5wpPDQPxvs9ro5mQ+kRD8dSiXfi9QsOyOjl
8XZDbhKWPT286eoZnjvDLKlH/IVYmVDLdFd9Yg8Z9Ojcziat9SZHG9X3QhLSrh/gQfjL3G3AJN8P
HrJSz3L5spRAr61VwL97aKp7WiX9Dy8pA6ddU4tWYYHWIvhrgHWe37B2SV8lWyJzm6gPCY9iyXC1
ik0Llg6pS+5k/5YbkcA92sTMhoMrLXQpt8uTKgY27pOBPAP5IxGuBptiW5bzdHg8T6h/BgEbRMeD
do5e3DPxtv7O4XGPC0Pya0+vF7mPr92jEf6VWVOgaR5WR1IcLQN3+87256h7CLzvrS1K7179Mnd8
RwZauhgoLrlo1TWSPxOgsJQsTA6i5ktQqTkqtHuUFfIzFzERrBx8agb4w56y59zoNf53meXkLZC/
qTmatDUKycfVXKI9j1Y7PJVrYra2hNlr50sjj73ruli3uRqNzoEwAAfopUynXvn9ftvr47ZgT1lM
7Gh0AXwneEW+wWj5BpXyc8mF9b6+kAeIiNxLoewHK1yuQLaK/iaSouHmV4DcZ9kU8W8mLS5jI9yb
zrdxEq0mh/AHc1r8Be0Z0F68qYrpHLMMXjlEF0fqimBBpI+oWdA8tgAmiXIAat8EDIeSiWOU47Rz
NxZ3gCIQciF04zJFs+qzVL1slwxg3M0WQFh+s98bNhm3Tr568ho4AVhmfd8Uu08MvtvRJ8OPkcnB
BqAvY1tmSbuIxUOOyBaxnyk+dzHpUldNxQc6z87U75r6XtD2I7nxNCELpVxXGlSqgNUVzZIOMY9X
n1TUl8PDjoTyI330x69ukHd73zdJ1lK9g/e70ZXcpxuh2Pe9VwIG4gRL9tJHH+qr+BvrgxAB2Rcw
b+deAuR+yTSp+wrvUlZjj3NatkvzzjBI/kqhN2J+uHFawsNKFZIMWNctGNc38Qi2OHtYQOpiu4kA
JwOr9mx8VEzsr6yDCiE6XqxEF2FMGwcNN8oeFavFosaek5sS8j4cnH6hJDJeNN5LvOcwkuz+kZVp
vgVFRDz7IY1IAoXIZLsTO47RXcCSA4hYjBiAC5giazQcWWuXjIIYHxQskay+ZikW8uTxo8oG4OnU
LBKopsRX/8VUhBKbwy2nwf1qljO+GX/mk3lZvFFx4oGofSIXMpSCfWRTTRZcytJrEcGa3hTjUrkh
gXADVQMeG29xdBIDyK60ILUlpYopl1oem47svfFVObZFpu2A/YxL9oJsG4m/mdOCS/aZ+P4RRW30
5NpLqn6ZAdC7K9YlhAOK2k+d+DSuNbn+IaG+aVeFgMsoIPXHEJ/2tFt6BzBOCwbUEjYRnTM24LAk
04MKi4A0q5b0geJUOsycrGeGv8XiJlSUQq2I0wrbQrRwYqJGFVBcPMeC8Jh2JyX5v21+oltqR/E4
4yT2fl5ZQYq4b5lr5EmGQOs9AncpMwncz6nwneM/pwGcGa+zTdgquwZnvDc5sfYi0Dz0DTBMD7C7
qVc3HZIhuNNDT17aaY6oDsxDVnchvA3r+1+dKALPvXwYjEp/WPdUth/bYiOqZBARReYl2++FMSlU
Uhu0qIrB6TskWGeNg07pXJunVQnTrfRnsNiTStKSloT1X3snSJ/h9mPbdTZGxEPo49gElvfN/Xwt
uJH+1T8ItTE9hv6/fzLsGGPJ6SbHhUgXQwUxlAqRU8FbLYRfaf3vO6jQP3c7eDGlNEb+WdNFG2jU
zH6TvZrEwWAHA6KGsWeHFMoWpeh7NJIwzHPx40e1yH8YYJl9VbIh5E04Ytuu5+05puxtvpYuS+6+
6DFmGuP6F3HkMjSt5hguOS9XiqBqheHwyuZkwd64dKG9sfnzfOugN9sqt5vQ5pg5BIlJboGwJX0q
SO2Pgq3asUiuPEtD6DjtSkzDVeonEXvQo6emNjFbleEpfOwMIH5i+66hVZ1ka8HnT/norOYkpIE5
G+YPr9DEw0i+KCHYgUvGtb/J23ATfXRfzEPZww4Fd1FzZH9cBR2IUPF8IyBT2Iro18EobRFZ4/sw
pfuKaxeF71zzogKePjL+EwdwlF5vyRhe3JO48Cfz0FnMp9+U7WxcVJRe/AKG4i1esvz6SvpnWkXH
mexmsrfwhhgwO/Y/KHXHsqzEmm5Xp3wgvQb0GCTyZBR5OcmverIs11tsXcKIT0Xcmr4SvFLhJzmm
qgpxLxKBU5EaKEg4WyzvyATDqDRv0qcn98T65euqc9GWKiSY9sZyICspG0I4pzK6ecG4yD77UzIC
7S6qpw6dDQSAPwbvS0zMXNxRgG+UGp0BnqcLpF/PFEzpik1GCeWWXLKRlf4mqHduvZhYGT2oz+ao
jPL9/OOGvg+qNHqhFZCwNS9FEmrSBtmVvGwzfPFrjoSNioKL++t1RMeJkFHJFPUIfMNS97LOxg3k
mK0+S1pQhihxqYH2P6ALEzBsxO8yTj05dD+0UlCH/b7Yi993e880WvPzBQ1XgLEbmQg9RHqYAlfY
aZFGZhU5utsQJhROPqYHA5hiWB85gVmqsZoRl+3WPoic+qMftXiyLp6Oxx9QlZUV4zBzePwS89HO
YNu6sTC7VGhQ93qdh5JqoBmSd3ZI5S9XbS+0AT8eO9frTSGEkEY13XUgmjx0mNndj3g39D4gmzGI
Wx5s9khL6/emdHvBvEKzl+Iasu+//z5S+R8ow01Ds8akhCvUK4RST5n7lQlGVxYzfF64EVdOge1i
Qps4xTTrr0Z5AoVigC63FxljmvUWeYrBcPOXMbzTT9+yq1E2TXHypKkJEKA+Ql7wE9Cv5cx/9RBt
3743c8Jm6JGsQijaM16UQ0Rdb7ehf0PqVPO8LuvhvR+zK5KmEgoHrKUdILjrpHGwHwqaUG24Yij/
ZJvI52J97ZMf+tHyjLi60TKBM6R3/P0a7/GMNXoe2lA78B83S9zS7ZYNpMdl8bOLnMIyzn5Mu7b1
jd+I/0gqHwvwWNyLScZB7rZCapNh0wcyaHgUz2TO1sjkH/AnFjWTPGFzDR7QWEmsReA03+p9ymAr
L7tFgbGeF4aoAtTlJuwE2neCJrFCm+u9XCk5Ql0qrNVSE/MECY3pka9h7jZWjvfi1tJuXxAmwdCg
VFmh88o9q9S4tvF0aFEXQ2tsFQXPVykcJTRKCxz5BAJy+6eYBDQX0HKO6tJs9V8wbI/+C49kCFxK
/Zc8l2quyPAehBUOqSg2rnX5PLO+Su4rxn8ESA9Dp/ZqrABPSG75Cv4B1ZzANabxH7pP0sHQWkCH
Y4m6hl0cp9PqZFU2Qkh7miomkRy1gtFidomnGPLCbpuECH6zxa5Pe+GQDnFWz2vvuycsXDCcTJ5/
YPhtRrqF04KiGISg1C90aqcAx53q6peIV6XXzOctI4k7i4E2IUfWqf+HiQzT4h2WLNuEUYZrv9yp
bpSUR0CDSBBdh0wqu9ePBea0wLx+NAhvKwizQRl9nRM7OB9ACRQyCLT2OU/pATqEfEig/tGZ0gvJ
k6DhUwbcP1IzgkuXOiI3SmOaHmCQ9g2w81ne8QYWtniIssPvvVO7r4gSP7F4pCcYcY2HSxQweqoq
IlMt4lfXsjb3i0eA2hIsq//yVVXvB+htNIpiQ5pWPR+k5vsQiw6NZCkhe9xR4kZ/b3HT6WOFLIeE
fgABsoS1cxQLT+AKptDWSvtqMkILegxxzjKCbS+SUjZCViev/XcyBepzVQ6816W9WJ3ND2XIk3F8
lgoSilFvuv8GVb39F5gtbf08H2D3fLvPnljJkhxifduXuA2tT4g+gJb7JqvPbymHchslo10xLlHM
QaMIV3MEgDiX7XC0Xid+9DWVHh3ix5i6TSS0a6eT8Y4wC1XDjz8nWRuc1C6CLmf/vdDEuwy/aTeJ
NXbMqHaLJGtrgRIOXP1QcmvL0gG4QsS+BDBn3mY4pkS3l2tzP/efJTl9gUUmLTM1BfxwpacOHikM
zxY8pu8phFdc5Msw0WvMBCz89RUHmxp2N8iiSMCEga4fjI/z+5q0tSEkkbnt2/pg54uaaqVxGBXH
LKEe8zoi19/CmfOVAeaYrk36fAM0qU3aMKR4zR7cPnyutRpkoeBvCmop6ESZWLMwtzExm1fiSofS
Ish2fIvXyKrHCZRiBEv0xy3dFSprf6Y8T7v4gqcX+7p7D9hNQ5XJNrTU65cAwHjJSbzJKmVeK6CS
dpBJIAIDCw9jL2VtsXgjPyOfPldzrkAfnyzrVgq0C9XDA+Jl5/nm13Gt1qDN15s1sDYzSDFnTQIh
v4BObeNixknDvPvwdM0vQwFHDNk3q/qQ/vdo3e4oJYg5TpQ2M+OrWBSHwu5VfmjBhyTzSTNG/DYD
oogkJCbQydVb8vN3Wq725iiSnyuZ0iY5tEmm+TXxLRAoXawfgP3+jYq5fEDExqQKmzsI/HBUa6xc
ROaYlhVfwnQznyCQY5zfXy1x6IFqP1unDFSFFbhCcDXPjMqyQWFQR1eYfd7DtCqQw9cJ7niRd4Ca
WPbImsryaFW/ErLUEgwE1oUN8mUY//4k6XttH09MM6hPW/nYCtaOUreY4OTH19e2LrmCU4xNIKLb
JSL86qLRhyJTKd3Q5NHjnFSYtA4d/5ZyJ12hzqXx982cMqXsYL4UlfBD+Upq+jCGSvXa/rNborDJ
M01a1W344w2mzn7rb2AkuQ/pulNVmPEwHn2FZ1fMSDpcvICb94viNOR7MxVfJibA2lvT3iRJaaXi
Ziz1SNsC/JRQkcy0I5bCGUr51OF9078TyjrFIImcfMVC9ts1XOa7jeeg3twaNb9JVOcy9qzySE6k
3Pqx5s07pVnnOUFi1tJmqcerFdNiFJzqCa9H9/q5+msxN75lr1mMV+rthhnIqca5bdWb8myursKf
zSX2cb23iZZm+0IArvTwCgZXGljErJN0TMM6ywkwKWZQUF4u22mIq6DMy994sI6SoHOoMdd5J6L+
pcPLIhJrIkUTuwzqMN0B8jd5Jp1WD1gZ1xleMZ5yMN/+BCg46UO44gQOCfqpsM6wPsWcOf5ZLvEL
cLGJ+qwvCWEgh0LDe30mlyJKUEsnupwZYJ8dIIw0Ayxrs30RT3eRF5g6Z3nVSN3xY7syHwYrJW4k
FoJJ9PUOW88AsDTUPvjSnWcpIjI3hMUZuHnJfKCaOGSa9LiPi6lcuFVPUbrZRVwcRG/ibyCn1aYn
OebhDSFQDCWSZhlqa5x3vZ3dGiApoi4teefnKi61SxL4z2ZckwCxeXot/Q8a76h9K7CHGvl7nIg5
CHJHr8yR19CS5zwKXeZWH53OujuLlK1YpGioXVRg1Ta79EGrBTFOiyCrwM/fMqEVF5bo6vH+lf6J
SpEBIM7F8pE+VALoRtHfzOEDXK+bhqUyNLN2BsisDG5iPeBjoNLV6XYUHf1SRZiABzaKWP/DN89H
qyRdWp5fGWTOVkAJAnbYkceKtNppYX05Obp0T4cGk9zNxgyRpJAD5iptwsNn+8n3UeigkJXo2XzC
+sMj4McRUEelfgg9WzDJP2z23fsxt9EZJcI7O8M4h0NaBivgTSFjpszsIOPLyxiYL36orKZcriZt
WLc/Zhzf/qk/MxBNRY2qBCXPuYvOGpmmtSdTv5C/5pdMOGEHxMWmvf5935Xu9VS4dXOJjMKrjwGW
kcGtfESfibXgMK577CL3y5vWOKGsyfzxvQN0hOsz9Vb2C7ToYi5fNnjLU6tjJdMKg9Jk17iU6Ogm
1l79kYhnoxapuv+A+Lme5vXrPzKBsBACWLi49b0nU4haJQE9fvjBcxhv0/+rVGbfoP1PYt417VwU
f3edXI40Njh9IXQ9lN4KwR2NdS3PTR7PUfs9nF910CrgSqbqHhvgeitlRnbZs8E/iE9V8h7uhsH2
BxLi1pnPRfaaRoMrt9DCqO/Mb/4ikMJqJPFIOAusdsfR4SD2FO+wDQW0X7yv9/+d5TxAC4ZmEtSI
/RxK2yddh7VH9NJ4BaEqw48eyjxz9twYcDv2ihjzOSf6befT/0ZBMN7hhSQXvV+A9du/nGnYhEhh
skbI7SJLTZWXYs2s+Pi4Hw+HF9Cag9yvknod6TJkQ1IHxN8ULme0hi/yB9VOWWWvfR/FcXccwyFj
s3g8QHa5aScJ3z4JaTgeyvk2Qk7VrBWKfkemcUWumUJrDSEDMkyBvbiNZ23YPMgHvnw/TCIAWtpc
c79NCTZhwV2prN4sVOJ2oWzuuxcNFD7JCXWD+SBnoOUKZ5K5VdnvIK9B47meCs8bbOvxvbtMu2Rq
A3xpzG3nFPw3d8oGeiXm+lQrEl8w9X7A/XxId/h49gZ5MGx3Z3Fu7gT7pYLd2/68UJ3Q0FIjaIHc
Wpjb1J3OZ+ZhUVl64rzEAmZxgQni4CZ6WrwusKxL6fiRN/ok7y6PAdJxgcvhDEfnVYkIEagvh6Ql
1Np2N82+S2BIkeZPoeVuUoFZPRZmXd8IOrCaeYcJBEpsKUjERixg+Efj95sM9iGKimBuk33eY8tY
ZjcjWWbdPQ0HPZfOFIb9+/N2mKH6kIkH/cCyupPakYGUfrCUELx315Da8PzkYAXaOXXRuqjkw0UA
P9G2hsnG+bZEbUS5LD7d0IGIEDTrC/nb8e2S4MglOIznFxLqEQ3mbsXkudc/pUyYl3x7tec8hXk6
W4cU/FXBhdRM6aO+yrF4rjyLd6OUS48f89blglaG6A00NeBsPaYZjL2LlTVnq5stu7/dG8o8cb6L
EoOrWqOQLM0sGx1DDJoCcCQixHp5ZImp1G4PbAWmT2Y7iRC22G/agUIHb+nsJsq87HeoAYjQ65Gy
1/mnnVFTQ4lEhnh0KVJ2ShJrd8NjQ7AbaYSQVzBVv1yvhq0uW0j56QE3rZnlOJW41qs0Ifty0cdZ
lEZDcSV2nqYKPUQq27zO+CY1BzWZxsGGSyDwNxGVvhT+dQmkb815F+QuWKtIMrXbEbgzyNKkBwQD
nSW5pqWlnlpwRpzhIa4AVFeU5lBRAUm+RWTxvuCWX0G1rrhI6eoZKhCvJf8P12qNwfOHPHwqfj44
FgMAsVUWZEN+X3e7SQpyqMUS9xfgI/iRSlu6ykB+r/QIPmNK8jTtYrWkFJDIqEBq5ICpOldNy67g
gV4Fa2jWb4g1hb3qVQsmbF0kFYDV7xyWpGZT1jAtI1ANhUWLDMsrl/aa16sRRTKbS5cCJ8MX7iRl
LzgWSGt3nkAzu0Qxi4yu7u4bbnX2vhnxPP8F4DZkgcC/O3teJ498BB9y+bJIJdUiFyycy66wBG+z
bg9he3h8E6lqzj1s2LVzoI1fcmi3dGNC1SJZXSZo+7vbHWe5SIOtNr09ItA8bFmsKkG8xIX5mTdh
TNIgAQD5Ha6wuqNQLvBy8S4DZcfToczgd76xc891hf8swFimQWKY1u1ifehBruhXlvlZgd02J/Ov
lhc+gtvqBlsh858OCwu1Z/7eS03w1Ejp1cHdr/AUsbXbgkGjuGXpe2uU0uLvQz5eQjpOQosTdLcD
cG0PxZFD7C48O2PfVrRAfbfJz+AcLy+s1f33DUYMpXF87EMM4Xhj6Yfdt3tqRI1s3EDXEqOvPrfe
JU0GcjdsBJ7EN2MJsmGCBd+4AxYnvmF9Qu8TvQ6mzOCPfJZGyMmZi5zYgNhA0c6b8uepzQ7/Ffka
0CUQA9xyp39lx/1iNx0tDVTqMqsEaYLna7IdDO35y8Elwm9e4oQJhpOcYzENsC0fLS4ipO6kuxWg
9kzr1yJfqeQ5HyuE29Urag8YXiLbPlU47fn7p4qjxyBZCYuCC4qCvx8de6OhQ5tPW53IoApxsKJp
427WOOWpxZmJfxoYVcv6QTIyR4o2DhhgVjd+bFsmxpb1fe/nDd+74vXd49MZS8gzVgbOHrNHEnm9
K/GchshqDuSC7JzGRjWB5124XWrvMz1XjaXvysqNWpMSkESTaRFEB6q/5+J2JpZ00EwvqaOPI699
qMV25A26sHXQN6vxcGTZ/cUCytFiJeXLfqAlCixP5ZYv64YYC9Niu4201IanYCG/pfqFKiOO7gi7
Rv8YrOKEhyLoQsCdyKJ2qD91ZlCBNpfOJehpUSyqBh/9PcI47wCTDX5YqDb02q93TDDFuDJFF3bo
aW/Lo+LCndWxIwwsLeVB9NQ8Tmh9s5Xt0TYCOe5Gfd7ZWvjPBDK/xwkOtvN+KLTllrnNicWkLYDZ
geIMcxwT763BBQMsBVa5MAndLqtxcSrVfI/0pXlItgsDlpoACrUTY7oIycfpEY6iV7ElAseBIHp7
bUr/fE9Svr710A6FTA4TiVUYvYXWZxFvGiCIJOxzzwoAjxEBDUrn3lhSK2vZEuoMEkCZSjjfOs3L
95zbtJnh27Jg06IiPvBNLIGrDtCW8bWa0h7YHw3DMzhhSkIxhrsw1YoBwiloDGc2UAVFUt4GHoRA
LqATvxFGOWpHa8zgW5wuAhB2Dv8W/kwfaAGu03SHlKO78N9oymdg4FSfHpIQPm24eCMxLAVlnf8R
58ioZAKN/0XT0Z1LwIqdhLCDU2gYLCQ8HP2zTCaDKavwI7hY3aemvEhBs+DBY21k0/1DrOgRV2Uu
4rb0h11fWVwV9cuu9syH8PNG341/m0WcrVO5AqLhhTx5Mo8tNw81+a/v5WPNZMEYgnsDzmvKWHYz
g8obFSmKMyPtZJc/ZRneZ9TSBMUHqf7thwbZrOMZTMpN51Q+SzHT3od149xV4VxAzujp9UfVTb5R
KSNc/4EuwONsGbEyXwa323JcFenSaJRNVLIHXwtb4b5FbILaOA41BX6gY3gWyzdz+Vb/vh+XT6Ic
3QI9qKz0s1s9PzSeULa+JojLbD0Hsn3G6BZsjjt2rM1F4O7pOeE6F823voJWn8d0Z6LdlEKY8ynJ
Hok1TF5ymOUXdpH/XsOQSU5foEI0i0rWxfSSvUKdNqJnun21fFiGi3lSz3Ak2SomoUFzj9FRoney
M62EABx+b3kHqrfx6BohxxjXo3sTyvDaOJvJ1KDFHyvFxmUilw1vw19W+TLIn+0PfU9fzMBTV/hn
FgHdJPFnz2CAuc+dBWKDHiDWwE8vTrzs9REmW9K3Ms1PtQ2gyJkzW+WsnCpqteyqJd6coB4Bfto6
AKSfa0R1W2uMmMz/tVsPwYhhKgRxh0GA4luYONDP7rx9ofq7EWAaIb89cM3L6We6hT4xxfLkfVo6
ZtfvFQ81AxpdtqVtclLx+6uMaAN00HlMtTHjtfmqwyiDUsE/AvZnfcZUtrcNvMAEWmPTK2GfZLgl
+Qa6nFaxCpc2cANNaMOi82dBjJfVDpYBellJdcna09Z0ylhGDkKgZcjdfJM1JPQfGY43lSXeVdO9
awxVHE2HtIVljcbrPTISnpGE29P+ZHSfSYQz4SvPDol4qSbYvrGix5H9FXSn1OdTYk30v0YHGB9g
DOV8pBGuaZj5flNIk7RsKy+yFfrmbjLwUPiySSJ9o6uv/YZoe9jHQ+n61raAtzJpu/Jg9nghBsyF
twUtpnRLg6l8vU0xWVOn9R4oS8BHSyVFokCGFei4B27UuD1Nb8bXeor8kgdbrivCKaDS93h4MEc2
2L2MrzUHouEwQmw3UvSW0qb9rq37ZYxcTuGc/s07sBoBI+ih1Hxh5ntdw5wiXqfJPPJQh/ceMx7S
+7jE+dCtFiQQTZVDUzrQIp3hcQ29CTIf94DSgTmKELc6i41rW/wB9hFmo3GzuK0DQrOcPI6JDlJr
OnOLLtos/53L3keP6Yu8mg6KHKqVPsTQ6hH1Vm2+JqoHCAu65ebdO0SMM9js8aB6YUAroowh8Nty
PZDk9gjPvy5yAL9Sycmf/V5XFdirJKhshExIVDA5aQkckit7xrXK7mkZbgGdAF9S6vrgBI5Fnx97
fjsga7AS1j9CJeObqSIMueyQ5ii9Uqt/G56nzuyX/BjBkGNdxKOaZpYcTPFIllfQ/yKGCj+ChQSC
sLIZ+oNe93f30spVLXwUcoXWSTiCEhGMEteC6Mh8dUv5e01aS4AQ0qlEH1w+mhYzbgpgGsR33Jxl
qsqplI9vckGoBy+SEW0XAqF/xq0TutaE+5wDR0Fe1q3/W8s9T0eU9XaFlccnmG+TE1PBwNZ2jrAu
nh0BSOjtHygdXIuqaEBAV/7obABoSztz8ubiJ0mJ/WDLcspSt7ZMtGKwO+hcIOk7PppTdoXJm9s8
mps4j2felB5aPkggxk+UbafaVzhFhTiMs+NqZp9bzWwhILweJ5Z6C2exPzNLj/Q2dcEIJPPVecra
2HmVGlbGd5DWPih/4CBVlsGFHCERiOd4nS5xZYtv/LDXpKojCOnbzVrz3lEz0jeC/Oi0Qu0OIJcR
lmhIf/rc2TI0ORfQIf1zp2ndFcEz23ZrPEoLnrIBrIOft+wa3BPnee/4sLLlUUDpeBnJ684zThTf
kRO7tKU1vQkIuFztg2Kkf8FcA2VYoU75ci86mq4e/hhFoa4Z13Wlb9CdJvzxWZaFt+NproOXhYys
sn3GzLbKaajRfYLT8qj/auxmXIx61fDDhVKIFhIjb4hQ9qkf2LWmcwHUQrmiJRJWR14XV0PYj0zM
9T0ZrnuQxQzyefrW11M+zCSoKNlkGUpAfBpebVUuFav0h2gRjlBykF0GbmbeXLqWR7RqBfE4cHJq
V+DnyDfgeN1S3VU0Mxt3Nxlcp13CIRlZxSqyv7nEGw0GTyQfYv4mqLs0hfdmSdfQAKGCgzLHVJ1G
4JWVX444Yz46JtP6tTa8q7cpFh9ZSeyQhwqbEhxleLn2EGFUnJC4uHnSJQAWOC5wIqTcmPVJCRGm
2iuKuhWUc+SIN7N2m9q1XuV7kZll/LoBTMrRwiDZ1jLru7+6T+BbRwk9oJDkvIQ2hJWz7WXaIrxJ
fQL7LRixJA71apvoJPYVpMT2SlQCk4G/yTdVX17DytInvJl3mq13TTzufOeeexAsWgfRi1eTE7in
oVr8mmE8z14NNvkT3NY06TU4YTnxMn7HN8Ue5HzxxyOxP9uXHWVlSdBL9bY8CerW56TP7v9QEDhe
PuQ6FpHveOOdmsBi6KdJ04zVPiyg8pZCftDFoKOHldRNNonCgEXZjAQ6rRfiY/WQFQNZ0QL/2RFJ
sAi8gM5PlLv1whqCRi/AAQLQWBphVJQdwEiaA3TweOQXQuv99oZHPAVMrwu3+PCsPFDh6+s5ENTc
hCVjivAFMAkNMOtq8uS4rHRTgWala2OfhIc1wEt4SMuAVj6fVca+kKEU9OvnfMyXquIO+T4MZo6Y
zr8Izffbr/s/RSVehJxPNJiHi5/9ZMMeJALX6wkFFLJ271GMGyZjIRhe5FA753ja9WKgaclrPRIs
21H6ZE1RNeAVCk67P3PYQ/q+hwMrA0Pa5AK3M6SeFWXb8Tz5CCcFVNSuVRsMXglwQVqyTyyk+4u2
w7JOLdOT+JvnezKWozdD5hvgYTaik8Dl637QRvSlNMzIEN7H7cRYTHltQ69Q1Z9jjspUB4L+57Go
EKxWaKkKWx+823WUWmwC1Q8dJNv5Q2Ps1lQJxBXtg3sJGM+n3vst5Og13GFyUQ8icb4pl7uVKbW5
3Vw3ve+1Moc3qzwpOltRMXthEUevMxUkbNBhvLx4EMVLusNWX8e++spKPF5OkbN2CP9da2rs5uBj
Yg/jOHjgpyMq7bcldEraP4CPcf3FErKWmPwr1ZRXb+n71DOK6/vqSlR3tZ1cxo4K8fW8n6kb5tzw
z69IOCyTf3hHa+YmgOIzPmHudsNEuMq3f3zC1u61fDv5moZmw5sbC/9VtSX8GQ6w18YusYiGG3nB
PFCL9rvAebAWSrUVb5HccHr8ev1SVYLcMnwHhuZaysO7TS5uJgiq8oWktqSSU2Gq/8AcfMvmh9po
rFSuIwWtPDCSMhiB/0qhJrocfEZV/30aDmZKOiwykVLcuu238FMq7WoVVcFj8OzrHhCRUkBbhRoJ
wpJyLtSilnEkMuLsDBDx5dkNWxuua0K2p5YnBA70E7IaChwHvCUNzr4aALALC7Ry9f/6+Zter4+c
3ROVlYVEcGy1guB+Rsk6DF5zZvqkdqgo/4iWrP2eXUtTPOnwrMtRD37kx4EJGa2kRo7kSsxpVCCz
kA6anJ/TaZ8T8Z2QwKuS7MandAUHhDc690cPD6hDfk2n2/c0qhiWjtZZORop6vxc+VTN9HEUpVB3
CPmqUn5go99Pv5a5g2xyj34hex2a0cbyRjXp7qpDqD9ernpkQSPqRN49EGSk4AZD0jlaWynMg9MQ
PJM88wgcmZ5r69WftviE0oFoh/ewsuRwikGv6jmJP7Mx+ICISOGEpVHJAXGlcVCHKDypo0m/az0f
+KFB/SqnCoH602b7diCzuDfDADPr0wbuok6sP7oxaWI3qeWhYDjRoixvxNUFF72lToqzVB7IxzNZ
xfHm1W3uQtHKsZlIPoxRp7rNb7dxi4BRjlCLNexrtoB85oGTLfgWkHz5GiXitr5u+gHyemEoE7pa
1qTkUh7sTKCH7mqiKOSFeD0vp788xlnK+NiBOaSllYlhP+4odxxP2yXvj6a30cpVst69H14STnyK
3VVqJLei9Q/7U5K72MiIQr+HLjd0SM8iKKnnjh2Fw+gZWI/cGM7ItAw3snK6Eg5S3R5Ylf8Vz3tB
LOwKxMaLzuD5gmhmCAsTJ5/Z52D6BlzhUnXjvHPgvn8dDgBp61fHg89tjecJWAXALRpYuXAno8uh
qkkkvtXYUfM+tAYy3a7iyBwgDkhVAlgh6yfi1ZDyj83nxfIEcd6Ty+xxqbrZwSMyNMwB5ib3ws3V
SYP91wv+H2UoPBf30319IzkAJjlbD5afNVgiY9un9Vt8Efo0Ota2Fy3zGW6B+pGJZ38zTwp26DRU
mwuOTKibiR+Im5mqQguNQ3fxfpJcaRiWmg4LtSJuao9P2TUWDE7mr0Lty/1zCPPlTFTGz3Q8ce1G
8VGG8AG5LDq8Ff2CVQMgWjQTjFO9N7C4QU4RB7KT56lVhimpRq19p46NwwUVhJtbcAO1CRBurawm
ov6wVUcwEUAqHhciPk6p3twwx0HZEVZ+Y3VKH6+rjRSmFHw6oZNjM+a/FA5QPtQaJ+jrp8GF05ZW
cqll5q5QgHgLqTNV5Rq+12csbBksaaR0PDSUWJIRbSdpojlqmQcKWsIIvsMQiBILLDxqdK9x/Uke
EuQfuEEBbmPm9otcXGjrMd8bheSuTIs8KmldISihsNWnh7jPTzgTTQtYy9r6o3uYId8MVXwiddxZ
2nao0+xNCZSDipRhz3Nvo+2absTjOiievaNEGdPurhiNdnohXMhunQn1pHYuj23sEPYAEKuVSagf
xxrRF12GCvw81PB0e4jzpkyJlhWxicP00tjlwH1TSSs1zu3qVR+u7iHzKZw5kOvHuH7aP2GlcO8a
rMCSmZYUjOJc4Fgp4lOwS81B9MEcBkRx9+Bt+0cN3l87WdA7dw3p1phyiv3z+W6ISqEEvBPRu7rc
nVeSh7QZJ0z9V9n75VwpFPpeY/IMwwG9q8wu3xQdY7606LhpLHtko9x+z02Hc8dJ1O6jOJyONQUK
+hNiqIM+UtYnkU3XIU864qVcFJUOoQWjArjJ3rcT5MFGwpTjbooCJvVBGg9XZmci6xK0ASnCgjqd
a4ToMH2HW4WmL7mPGsYDNs11syR3l7fiXw53DGMebOX+/MgRjH8BAGY51jD8DDEf9NB7z+SoBLW/
E/hvoixQR/g+hrwn/AliLgg4HrVafdwnupphtVMffk9iQKLyX6/IMsIylczPOuxs2j2Rn59Yi/nL
6lo+0YrskdTIfBRDbY+hECJLEoNNSvkzcde+f9ISKLU6fUo6oADXVBN7TA8o4Yg2LjgvXw3LON6V
vQBeoJEbHFFAvP/g11bQGp3XoPLUWTRFsc1WjUfp0heeQvHxBmC4QBNH22kf7UkzeO4I1CLXFU1e
rojAF4tqaq/+1HOv+/qfjceg1Rm4UZ1y9bQ2mTn+TfVLi4scNy7H4+Y1exgFKMdVv28VnB85uKqk
tbKAQFswtYf2N5NRrhTPVrPaSLuepmhs0hGdawxZMhuFwWWR2QYicxwLi+HfqNGhyKc4uiAjYrST
lQupczd3x//4EsojaiHnIWr60h0bAut99DMYizO9s48vNrFqOyXMZ/Sm2GGURtqKMLk+t52PLhmV
R8TiHF8aZ/iADVaKGR0qYgM5CJq/qKJjZAO7zs8HDa9CaM8hR0pXegeyM0d69PqPqkeeNhHjULjX
7nDgvPNZORrnbzeJnzLBWrl63NJk0B2A8O+pY0fst7q6Vo8g8S+bR39El93aKprvZDuDlL+8EclE
Ggf89Ama8mmzc06ptIB76eOvKl1Saa4je4QioGpAt7LdHgiWTgVZACgRfzAZw8TQ+xSONykywnc5
3gWD+m9/YRiDKrmbgEaOx2cHFGZqz9n63pu4OsIglG1y9XQKG7xNjiVsvAZy/nO0WgVguBOV9Zbq
/1evg8q5md9bmITMcP2nBMKS/TyIWh2Tdw35xu7MWt7STkjnVHeFiEfDrqg/7xuU6yvtXdlC3G0p
sS5IchTkEG7LmoRPuKl8qyGsa8zRKs3iV7JG5RhXfkN8FosKPaImhXgyx5bmZDYnN3hbtS4aetc6
4yJ8yNCaU1ic6W+sVfLVAfMusr7WecOBSojVUNE8bcfaTXn7fXBXN8os32XSoMDgOmMmxAAGRdij
zGfMyfYEEk5Di4gxw3UfGa18emZc7CYOMWlgz5OvVmFRb4yXEm37bOR4LrhVoPindMMGJQr0QuyP
/CF7VjGzIUToBkHuBZz3dD0gxeozCGBDTOm4X96P53jY0mTEH5BxAVRyMcWmRa5C2fkM3gDn7y+/
14z+zEUROVKBKiEZ4bIFVJ1VBtfCqT5h5Kolwq7utO2R/xCWAt+ewEQhQdFrZYbWtKs2gyvq+UbZ
DS/Pfyif7RhLQ0esf1bflBgOfuUByDYye4orVuDrL9Q5mzEf1bw7aE40PgsME70PS9yG/tcCIQNT
waLounVmSKGx7X4iTMmpWyBDEdHet2tWQo3cmlf/acqi5iJMvYHx+GquTOnvXUMj6pikdOn6K3/u
P+FA497VDUm91ZvWF6OcrfKyk9MAJ8O/Q5I6YXTc+Uf5u7po+5aZ7TmhPuBHUtd4p0DhSGWX4bvC
LCvDA9twBpI+ptigaRHRWbV93k8ARE9cuVJ2B+UjbuoMopyjAS8L4fzBjdOX0WPTVp8CBnWc3hPb
wIV2F7Z4OCvbKz3oqJXtSFZet5eYLuStqu7/M8a+f52OUSOzG9lByD4sEMtyv6+jQWBWvB7Dxawd
pgLnQzVKtrKf4aXh/wyiLzCn4i8O0TckWv6pu3Wt7R2rZFNTODSOmRNxRaC1W1Xo526sQjiJ/bJP
7sQs/Fzyk81Udm2RqviTWq152m6bd4cYbmRUAU0oxNVHL7eM6hg/FlhfBW8TB8brZRPt1ggb6xUt
1n+cwPHrBb80GQBI2Aoa90iMGZLy/P0gixmRZfONXxUV2+XOM7OAt33LFv7Tez2Wbv8tPyf8z8eP
qeYTEPQfBVNsc6bKfq25Esu730Dn8QVS/5D2rZqMwFImjOdK9Mhl7EDhreSsHba/0ExJLvLXHns+
Nqeib6jI7Inbj2YiMEJeSZuvnI+zMQrFMgCkhxAiMSf+p6w7f5rbqseH/1qf6hrve0s5ZTu/O5hY
r36pG10vmzBpFTU5NMxuqw607QfYUXaSqdPUYd7oRZ16tUQpjHktSQAhGm/KlTqkZ/XIzDoLN5/k
1WVJWiexTRUGFW/Z2+ZPWcRQ1uDunaHcO7cjXe3Cm1v+NdT9dfVaadAfrk9tCzaXshaZNuVUkIqv
1QyZ7dpcIXV/OGKGj/kmslWozD5s1iFwK6bvXX9htezQEBKZDazaWCcuudnpuHmOgWwVumVoe2ED
5CbUrXTBsM/VVPXPFb44OsbvkaDjAJh6E+DdNPptMCxYXKgXBp4UabKGKbanUbxqLiuPQeZqUQ+E
SXyPR3Fms/XxNzLsFlz/zsKLQnbgAjgNvfuUHFOlKl522EdbLQsgwnztpDxxE7IcJ4EHkkG7+hJt
hG2vkqyYhwG/vO0dCroiMNefqflJdxdiFQMtHNq4sf/LGgfVlW7CliwJRjYTRlYjmedKXCV+/4V6
dG9lX9WavJPYRpL663yuEH3gAI1f+Rh5eStIZlOTZJ/Jbgt/PUCsemL1zJvzCnW8nIhxxz+1onNW
cgLOJbS/1hKx0laLMIL3oVqEG7B4xBzjGwtKv1yxr7nrP41j+6ydSCCE0TZLX+l+1qw7R8uM2XZA
piP0DgJhJCSP3MI8iT/7erxm4HVMIJa9pbqbGkld7VH97JSXqfkomhY9U06T1TCivS2HougBdQUm
YszaiCMTj3KpVW26mjATgVY+n+Y5ES+c7YUqozpVD66Rur/TmnP0yOI/dNE/P63wx25JHerEEgul
NQV/HELfpV+zHUtOno8un5KaMWIjtDWwdAcODRU3jAW+SRI1o/MyCKfGSMLcQRNDd2FUv7QosFMD
bsS/gnHIB8mbosIT9+aLQbWnhacmNLeAE/IGr4vArvKv4oS4sBSyPoEZLz5mMSfeNBZNzprlychR
0dDvniVyLCFRQdzGZflcDAK7baU/FBD6Aq/a7r8x/8cenKX0zCc4UjTNCdnrYqCYQ/M2dXOHLbfF
sD/HpQTOIMC00q/MstApAsvN+KWY2VkO0CTjUQGrnNPWOU3hK9spM205/t5bVjTspGHW0xpXXaiE
NuD9byrbvMNrxn7gv6XNXLhHjbwdpWz69d2soH174fwVnQER8qqfU3mcVWu59iuWE/3vZCHLR3SN
JymEiWKZVVXdzL6j2cqXsCRpfMKLkZe0lmLXcFcajLvSY45uwzYKUdub7JhUurcnXONyjOzg74h8
YtiGfAAojN8o3xJ8x3PhOVZqGPvJ0nFk5S6byjy+9orQT0lFyBIvZJuJGxCOm6R8zwG7VPwIPB7n
tW55TfoTw+Y/sGkSj7ltphPinvLwFjD+qocA8lfoNxYnFRXi/k9d5pxg14wNL7w7K1orNxddY9GF
xzhK0RnCF3Cs61kYCxFUjGdVUTi+BbQsAJ5o0BnHccyIwOsHAqbaG6zvak8v1Ly9gZZ/qY8c2cXE
b/65/pgTNXxsbPDx4Y9cgT8EMyoq7Fu3Q7+zOYPs4JDgR4E/RtUBlbaEA6GKUuV8osLdtMlMmDY9
V5Qcc99kefdioESoz2BKbKL2qBpmFtt1rRxcbzPsDnjbhaOIsnLieRaeiKLwvZ+/vuulb82yK4Ok
xA3xSEIQEm0i3CKcgonzMCvRzUmsg9YbKjwbI1SvfCMi2zmcW0ZY1WqrVt11wiPMEddJtrAytmeJ
9R3j7fs+nSraZ43oUksEQ8yEOEUa+0i3X92yYHtoRkF+wrA6m9eHNQEiheuQCuS8ZUJbh3uU8qw4
ikZNyiYpd+GuOwU/lj8JblAbsVwHMZn5PkI5OxdI82TK59QdX5elOGSyEQmXoDosRw1IUUYfcyp0
UTVzmh/ljOhZFUJ5nYHEDqnkS7MPy7FkdHNCL7M8vuq2/+d2gepso8ynuKNNSe8ohDVtqIPPz71+
9+8gOyLzIX6MtR7o6QPZo3dW8Z+A5s5QclL43vzo//HXQHqYOQLAkaigAwEgoDYZlzjDwvc9qXSD
xwOSwW2Bp94ODRNsB+oJSN3z0UyCUMo58NWPVvyhZZ3uLIXwY7Ircydp3A8OD2muIiXhOPxyYjWi
vH2WaUwVCbkbKb2lOAWfEfX4ZCkXHyLUcjX7e5cEKndqmZurKWtTR0mPOE14Nvp53s/m54GJlGxT
7EpM+nOpV4qjzBdlfKdK8eEgZG2jA14q4lF3hQKuWh1velqyDxZUm74rnLSU+dowW6WffrwmLsrY
Y+wDbgIBo+jE6kMe34NTUY/5esKd13heSHzN5EhCxfQOXfDj3+QWuFFfzBnhDdiP+OjTldWBrw6Q
PnhUHXH456DU1Tm3xDWgddU6pAAwExYixnjSglJXcPxwPDDdBg+MfIMvr+qPygXl3qyw4c4LXJVK
gbCilXso9R4t6VtfVdJbsxMz1zII3L5oVlcWvIAPCnFSM6tD0mMeCsv45yk2OBbR+f4JoVo22GV4
0mebPHPJc5hFQrGGyLpwR6LoLdsqtTLCW5Q2MY3N7RhP7W0K5n4Xb0cdtLAq/Fpxz182BxF45NG3
k5ThzawWv8PXrbXQdhZl4fQxMVwUflCTaWaHsJ5GBB0imAeUL0gOmxALq33WksNKlJWtVuDyGdxH
miTZkHn9FOmMvvcYYmkxxG6TI/2g5LE8ItLOi2y3o24gGJ9LhbErMQdy5ZJmC7qo4eFChosDM7IU
FjsYPRdNsPYbPFX9CCew1AF+quIONSB8o7iE9aIQgEs9lN8sNyH0WZuUUMlRPFb3EtDr9vN3iZHP
48+ZnFSf3buOGHbrkVbo6RK/iRFcfA5emaxrRslaPOOxVvOOQlopS/rmRX9pyWcTpCoF66GKwlM7
yWz33xBW0XSVHgVlTNfe3lahDY6BU73D8noLb/hVUDptOHWLipARL/KNeyImSDeY33+Z/KsAQNeT
RSMFwNm3ndBBmUzhOGt3UVZhXPtjzmtWsDDkyBu9oNHFHuoPx38hCWLoWyvqn+iZ8BhLmVlTXIeA
Xn+1MdrXDBD5X/lt6yWTujSKU9cMcZYen0mp1jA3C1xpscv4n6DUkAHMhluD71Wu0nkC7XBCzWJB
qI+lNF/pwYp7CpEhqVfwwaQ34VZfNkfNN5p+3L3CztOWFMHB6cJqX9V25UDXuUFvKJKA2uG039LY
o5y4PdEjLkB0U2tT4E1dSPn/oF1X6Ot3Ez7G6cEeKeCnfcLzbgl6OonUnhgu+HbY6oaQehxF2/V1
Vd6nSHXYWeUUkO4R5krv9k/udtx8763eT8qPwu1NDBpxqyBr3H5+6vygbq4POCtdJ9WohvuF2g5I
lFIduq48hBjax21oSaqX8aOZ5N4NFhAoxhMERhZn3C/gjLYNWwfXQZ3ohG3vwRKgtC/eRA4mdZnQ
kH1h/xwyknO0CxMBnz96C2M8Ic9FhK3ZNE8RyGMvustrRIVUTkazwT6F9fGizTlUzkLAJJzbYbBs
bKX6oQ2bTGUj9jwfGUIremXu3P1jBPK/lUY1OsAQ8lRJ+snydel4K67cbg6c5DCVzQnHVdXL63Ng
I5NKIb+SVgbGiKbTtLRRFGWO9Poo+DbeMASmFuYrxn0trJJrPTBSXgq14maHc1PPC8vfp9CyjtZR
hriAqwpzWZeD35h0GzOwI7a7tVjyx6p53Rq/tQV+PsapUsM8gV9EP+fki+iM3yT4crbybuMzqEjt
DW6LZviFc9u7KG1/NtP6dGNuOd5gqqVDcM/Be/YSbQTe/VveEuJpXybMhUb2ZVIVYXBpbWTSuc+y
jtsKqpCWaRRXohGLuiQemrOtC6eJ4nMGdmWNSBSd2rSUtVxdhjpIk+rZ+umjUm8y0MoxdzAmOXUc
uSdfFWdOk3fK/YqALhdaTO6vcGdOhyrdIelbJpRqpTrgL+ofKyf/MOmFgujMjb6gvOJtyVwVve9s
PPRk+kleGo+FgvESpHAbg1iJOC3PhQenrU1TqsiabH+vQvD+yQ9AfcF2xNeyw1qR3LalOzaJ0tKJ
XqCVJUvqjK3AMU3UE+ZcpsCnkL9VJxBs+ZtlzsZNFeN3vZuXy8+B19DGb9LNdl0xl9PqT9MTl200
iPFfBMER/BghHbyu2JR98Omu8LCOcwNJVZLKMn6dhdM7rnzBmv9lCHn5MWpDxtNxMtR9gWMgrLs/
IfGMzmANNCdJ4aTI88fWoyWTtxDpu9MC+2W7GHEKUSSwC8ZFLDiT4iSwwRJrNlt+RyhrOzeJ+b4F
IPFZYC5hgtXXjfzv+OasFTXsFeU5lIFb7m6yqFGzQnwKFiYEMtQGdpT4TzQLovVM5cxYwbxvUkZ6
uMDp6jVA30tTlbbZ5u7eZuuTjh5RWLX8rVnQM+7z7CoRGMziYhrT3xnzY07WhFw6VphwU6cWx2R0
XNE3fJmPgX9e91LLns8KIdiyL5RjVfZCKk/La818GEjaFn5nn/HogVn1e2OaaDKRkelfDU2ZKlHU
Kep2q6VY2RBvZ6BZn/3Qig1Oy6561Tjee49HlPiNIf+yv6Ia8uNNfs7ZF54IMLSSW7yy3levsN96
kkxpooApKP3YO5hnLFDcqiQQXHMbEmEjv2IsIRNlf3vmT4+w0u15EHrgOgsBhyCZCdzMD96if4+q
HRR9Y3hKrELAyXQ/i2o54TS3JaT1QtWtvAwcwzVRCuy2yfFWE1ZXVpFVJXmZmgQdPceJz3BkkxTR
+hIfSGoOXGMhS/smjJpiDXx+C0+Q7VrzhC+7QcI3syElb0K6IOxI1HQP/ESN5TiFQdaAeJZlmh3z
Z2aY8ETrnzzpnEk6Igvyq0VzdaXnWPv2IreHt7C6O+rpc8eRpRWuDweZZy1jw2XkGj6sMVF8ZPoF
i0NdhelmjbNLPG4IbMMyy58pv2ODixafyiCRXjxV6s/VIzBTeug3fyK1ZR3B/Zm4pJq6qasypglW
R+sJsG5d9yUwyKmgFWl982vj0ICr2O0KlqGX8raNzxUPBUWy+aODppMxPmfBqrAmLkmDPIhDTCq2
4G+i5heneGp79qc6f1B9vxPYNS2blaxLKBDXXbQ3J1lv0PvHla3GincZnQhZ3VG9eiRFIlJx5XmE
PGDGVLX9E59v8nCdO8xRWFl8DxlVg6OyUJeGoXW3AgtpHaXiZg10sJqAI0+LvZplcI+ndj5EdXrt
eStxZAHeN1f18uSY9CRdgroO/jOdt/5PPCv4GeOhB7dTlhUf3cAwFJwBS4F+zo4Z26+YjzsE0Ai/
tqPmx/lBOo6hafPPM5kZnqSsSYYBSBiWhClAeqo6c5rUjo38IW4uClk3Ec5M/J/+B3gDuJgy79OX
BJFA8COc4GTB6fBAf6D8COubOGXrUc4IDkb+Ptkqwq53JhFdxByRTrHzKBYVzKdi9zGv+Srs93/g
LF8auIoFZUzMn+tP3wKburFEQLwroYzq4JU3LF1HTXR+L0ZGsiW1iJNcBzKsJtgTZHbvvo6vFWTq
Z/HccDdmRUxTPMicZfwbaQRsg2JyPG4UZKiB0kHxyqw/3W1urLcMTNA9jGogFuC378CLP/bDqVxW
yoz0RlJLxKGsELjLzEl0pJYWaqrTw+ki9QxUOoi5KowDBn0JRcysthpdqu5xP8jIxS0Tyk5sLENg
8+EaWhbFkYmA61s32odAv1dJRwGuOq5Esz3+lAF+cgRNN/HVjxVSNwbc8c40+J5kC86k+fXsuqHX
9VB5GNldIm3hRMRwUNgnqKnGbKtu7bHmB01rBDLAUP5l7bRtB5i1ZFNuV/lsQ71jduNJ5E44W9eJ
822g3hoYEPTdowAUvSyqOdWHDWSXazB+5ht43teUYcCferKJMOJYQxpJB3y3WVvJm6fPHkxzf/5B
IoG+NZeRrAf7bqxGlfdddaUWwF3EY7qIRKaTQ8wPSXnyC42NNW+y0787keHmS7EW1K2BtB5K8c6V
Q4zLyWGve57qTP+FzRuP7vLSZ5zu/65nDAOoMw0xFe4JXQbg5+lZd4hvM7dqAHViDAql61fLV4wy
04UwGxtFvf+y+YNgjhLDxgmAMiLyk35a269bCEmtsXYSe3QoZT98l2plOlgbUYrkj8r+se81B0Df
OMGO4kLqrd9mU54qdKvx+WlRTQRXnxx3wY4WcVV0OZbJFXzeV0GCCmqujYq4TyvusgGhXGy66Ibj
f16hp0EZAc076CZMaumgXDTQUK1ykojQ+6JGipGDDZAMloxWVTOEzpesCKtiO7ACttrCjmx218UY
pOk1brcqs5jEn0DwhUtxfotQceYdE5TmZa5RE2rybOBt8+mVSj8FYfAxetVBz7+a9aJWUXSuxhyR
SUm3md9o8hCHz2WiBRVol6WYZp4AZrhmx2JJROuwO6xI9T3E0E/lQkiuBtPYl7m4M6G5zdSAooS2
xcOG+wm1N9EllVXK7iMERRiQxVQGLFJuSXDims0dUcfIYggIorbF+U9X1pR971iHKy7BVLsRFZzL
Q3S1FYP8w8ByU3HZPkrNiK1Tt0QqRIBaJ+xSbPZ0SwH6+wIJQyYbKcgSUhh0qfWrkYOTTojK6Rsd
GLckEVDZBICYAJSrWYW79o6RhLwBU+lWHWic3lqpGoB4Detu/I/Ld+om8sh6qKBz2QJSPN6taNdX
mkyHflE1YOBh5QJyNwTDDULj5+/D9aZ4t0iHrLMx2oxrbnwGMstFyUn1J12oB4+hQVh5EhG18nbw
b8k+ajLB0IhtRRZV89BOLqMx5y6DiikXNPNCZtpjgHypTHxEbMQhi9WlQ39TzkAwfGZZCq+89yrK
mCIJQOySe51GW9MWJH+7vyQk90Ph9purk1SLXjP1Ejh8jcd9U9+/oRlOxh3vpmeT4BS6ookyJjiX
+ChrV8foKyAA1B/x0i2WMQnTr4RORRCwzju5YZHVMX8Y9HjmUCTcouWQqVKG2wylrhZCGGO7OhVf
gTc4K/3g64v5HV6iM82CD4E4z8sc30oyaHzlYL9a2zVVhXOJg5Z+hLUpNcfIfAR58FIbhE/3GaCy
Jzg/VmmBZd/ikZ6WsjZ9obl0KnjwaKPZDVN5GvT6as2x5T7OXUg9PGdwfioXT8iqv8xPQRhUWF8u
KsVA9yXdIlSVo/fdY+XTk90c/wIGzpmKJLePZv5q2XYGn0bD2RS10ijZUWpToeHAyek3RZc36wYm
/F8Db2otQFgWJEVnuqDl7WtNGtBtipLM7D11l48M3c6H+p3Ys9dEKP4FdUHvJFY1OoD3CTkxpzRo
g41Zuhp5/xZowoQWswlA94RRMP1aESwoF1Bw5cJAnTzxK8ZXO26DUC1AJqJNxHhBrIk234kqyYIp
iLDrAU5qO8j3jDMQw75rrpu0pT3GuCJ7hJCwz7EQ5jBJpJfZWGTj6+CtWbq/HVP0FF+KfCEGUJha
vfkms8FuFF77sY4B5iclbcn+7W9JzdtNO7pCRalcmGBiQV4sFTh3fsqu5+bE6QYzaTEY6jKSGw8o
OQkHcyt9wBvBrIJ1b/Tkmurwv9KBf4+nggpDIBb7/+332r9yJrt52MJJ2pCyKodsIuQk9/Wb1g9U
zZpQWw2jEEdiHZ5mN6N+xD+0Q62/7wPQUKHIfcuWte9ju/Hwk6AJ2/r2WQgzpXKjsFMt6c2OIQ1W
bifpDtzYxGQiaAa4dpRt+piWiM9CI4HPxr5/BZTpEABDO6GGi80FAQYZhLsEKdigO875U0lxZDPz
orL8bG+/ssugw/SKUQdnwWGN80GYIs3iqGI1BUgnBPwXopgdmDxvXAHsLRP0aKj9Q1jEq8rIuT4P
zgyLqQmF7z1m3bY4vpVanevWzWWU5yo8nyiWtXB37tbXBlNNprK77z6pHvAhMEXJgL4HgcSMBnCK
U3L9H0DxQvRxzB3lERDVdMFo5g+mrWaLgXA+AKiGWnOjYWqL2dPxJE4WUL8A/PAAUeVcqQxOxX31
nmHyyAIHvPsq3UjE3GFH+bPcWIqbGhwPJ/DA3H30qEIr5Gp51Uhu1DeUPJk9gFSbOH9KjBOTwFpe
CLrCrneQzgOarIPOyml+C8DnFvQCh73s6oXbEVAB0WQi4iDEROzBDcrFJUlak6BnhJcEgLRmw+Z1
Kh3J6M/pwtvjFknP3oJqlrDp5nxHzPcYYLm9f8j+9v7XFYvZO6MSIubjpCszJm5GMT6O+oWt3FtW
DNz8+oQSt/WofNL8QONxT2CMinl0DmC2KCLcahXJ8W4r6ASTusp0M+OzJhAmtD7qEXhcHGZJ+Gov
NLQOVZISNeB2rgcUy/efeG+zhwyktJeQsbr7S9RcNjWOGAZF+R43pbDprNgu07dZsqvLBoWRN+Mi
Ri9CdAqzhYCq4plX368cBKyjC5miqA4uhUeNyxZOMfcV4Vk6+zXacygHPtpsBwOEqOdXyHAwUObI
tnr7SbvAtqK3OiAvg+roNZuKxogBKf7Hi6x/Anwm74TAIMPhTXk8Pw/6P8hEqSli8a3cCJZsSBD+
ViaOS4g1xzTwviT4aSD7PM4ajq6dbwwJxjaYcK4lmrqqBamiuNckF3x04mwI8GPxT3yKHq9ZzZpk
TVK8c4Va705159goO71Z9fYCF7A1BPnMw760fpRQ9bKdWba8alz1E9nw61HqbsjnQp4uMANkIviB
NTFYCvP7KHmyidZdM0kw/Cf3C8Ho02rSPim4Bf+01Ik3rfYJzbPkDqvW8v4DIc0aPQ5xy+XGiE51
3haGuFw2YtpC67DWt0UBgoc+B5zSPZ5UDIKxg92Cg3CBE3RQjTjLxTTu0gM7HGI9W4vyeb9Pr1Ip
z2u3IuInJ8RlX2RWdHRFyYt7EoWKsEJ6Nca2AKxmb/Wli99zTZSSTAgBZbPVEPsd03WFELMVXxrT
G4ve+QyDcxPKDx9h+2WZ/o8+xcy/KRowznS+/5vYJ+S15MPvo+fheb4t0Ciq4k9tJME30fjjS9o3
zBJAptpLKhqpXh2d6lyoZLKV3KsXHNfSCWoF0aVCTwVZ56Czfhlp7BWRI1whuZqSyEKm9xHtu9+D
JYUfT2kw9wlVjXr+W0c/bo2Q+OmHppN4RXNPts5AN+f44HAcWkRe+txI1M2JYhFuiI17ziU+OG7i
1uZKtGzoQsR5PdGlGo+Gb1uFhc1fVg0PRuIpzTAaCUKUhfGTB8n62tx8vjTPAGBlzcGIphjyBa3r
4u++SGuI+aMVgGFHBntJvQ8XMDQJTzs8FPxSKs8fFlm0HTmzYe6cxYIzRF71AvaV+Lf0RM1XsS4p
7HKLCKFybBAXEn50F3+mLAMW/lNvavW+DQ/cO6sV03ipoxFQsGpQEQ9KahSiMj5RfVlNphKWpkOZ
0l7tf4QQIxh0J4AgrwIQrfWC9CR7v/IQU1pFDnu4MhA8w1/qHWvzPJ/yaGd/bUwc+6/2Y2r8/bRA
OKCLVlrFAXRPh7YUqeDMp9Wz//mDB7Rnpf0agNsfcynLgpJiFsjHN3XuNzl3YoF6LM+oSN4iZbAR
/WaT8KjPj4v6B1fbj+G2qj/IYEnt3n1iEe1zePsEUipP0rS0gGbqqoSUxxeQJtb7uk2Fn29PbCHQ
AoDv40mrP4Bu6esEsxlBUIv4Mf5rkONlswnbW2XRVbaClDVLVBz9XzIMPcmZhyBzWpD/7Fgwsr4u
m2hDUifXTCfeI8rd2YUCJDOVFIlOdNX4ol+UShzFLy/O2GgJqusMQuNmWx2TI9l0HZZO7IwFVn/k
/oEl0pRihBPTVKBxtk266JP1PgaUGN11nx16mdihEQb+JADj6cWXzzDibFWRHTuVXIJRwRyBIUI7
4HFyKDTs1STMg0Z18kkJOAdYmhCH6pluGOydh9vJb2UFYmLxhExKQa6xoIYtkeqHsEKKxwLqP2hc
xy2VLzNulMNqaJw9m2KxcofCKfXGNxoZcpL6Jj5LtXll9rRbR6DJlM9UKTs1qwE3Kiy+4zUVxFbC
JNbT3NkbblQRCPXGhvXUYbHSrySbqwJfUSHfJMkhz9v+AgB4PqRN3D0p5HWd1XIagBPoyJX74wZs
WN2PbEF61gbdt1hBbfYJls9/F2tiX8P/sJdchu1vwzR2MYeegbtEGnlDbIQ84TELkhShsY5M+wff
lknR5XcX1wDUZKOS/j01uoD3ojvlGr5RC3JG1DW4EIsCCsWjMuERTb2is/z8fNzces9aDWQm2WpZ
pfuVFTgkcdlE6YVQqlPIwp/JYFpVeBUFknSHhVnjGw7TgkfuKC5b4YF/7uUCJRle29oFejGPGYBo
RZiymxveZwW90tkbK3MLbmzTmVwyLpaVsHnKHXAuJGKKIiGFilcVQeF17Vm4bwtC4doTO0rlK55I
gL6aQTSSltttK3QNvO72cq2bUmWNqyTZL250SP7kEoqRfT/248aZBYDETPmog4WOfJWWVdho7O98
h+0R9Qxe6C3IYv8uvDplgyCu7PTsrJCnwiQG1SvMCfe/OS0v5DKEJx2K6Q9MtTgsYWS7DOqC6/ly
NUWEoO2d6GdD/iMtzOR9eLLLExgs2BikQutfRTvWscf31ZMqwGO/TolPdeNuskLnqBiRd5MvTYxG
Qhsl++Mt02Go19V1VmNp+hmHMrSG89S2Q26/MZYrm4UPzHn0RPY3EmgOHrK6TUdBGWyFAlyJWAH/
OG2HxfQ/3T3VJuP2R/zAxkHcT3tKIdWp3OoedxHornITrRyIWtAv2UHe3EIsfou3x6wCWgpzeY6Z
/UUuMTjjn4dnfZ5gDEdjhmlCePxM0LEeqSd7c7HLaaf/t4jbdQ9KOg/Rq/82LxfWsfBsAbalLezp
IO4ZzhzEuqgmu859sEwJsG8nKl+aueK9tTfWJnsXXQrLuMAgWtKT4Biye3A346GDfbKg2sqFyRqt
4KDWxnqclUHiGrvr9LJrK3xpJkBxCma5XzTOtKo9ZjnfAqWKIGKLsa3vt+UDHayFAKZYftBzn0CO
lvpfd0lDO7JRsxfE7nXDDJxP5Sxys1h5HL5BjMWA43zxTUX7SGCuuD7KCx4YtErMk2tbF9SCq86K
HWWE876eoAzFIrIWWLXx1gEAzIKL3V52eRsZXticQKEL0cA0LLJN7S913PQxvdI3W0cB75ZyMQXZ
UTW2WMnoSKtLqrIfIXmUsYJm6ub3JeLuQOP/ST6EQPTnF0dLa+etpPq06gHwCh71fJV+pGfAEzA5
GTef4xU8KuaaTxqcOMtnQ3nXytEHfgYXRpEI6iD7BIjcYdggK6pFmLu03+WH4y/U2DhE/R0NkAB2
nbvAggg8ffPIq4VL6U7idIz5eo4KvZ1XYFytrXGEhCRWuN96J7yVuk2RaFTCL2CZA30jZyhfH1N5
IJzJSImMWIr0SnFOn2e/LEM10k4UFjJr+4UeEmI/nq1VGP3CIYdgXD+FSxngdO1Av56C0XKdVuNQ
CnqY8KYoxGlrXrwm1djeySWLrkCcyvPvvJSBnr2b1h5ktaE0P6D7njdBPS656vf0aPINiD0sRPMZ
Z+VvW2yCRva6EPJ3a0vFPZOqRMUfOib0p7F8BJIuXcJiSmycugoX9zS0okV8eiBmboHhR6fp9Zow
Rr40SS1CgiyLCHO1V6QWfntcqU6rzNg8DeOJK/qgQsSNq5b9kxBneKiJ6UBYLwL26N78NA+fv3Sp
ztEvqpFK3EILcK8XSU8yFPupnYnHfsRMhAETo8DC8oj/BPc8nJkzH2mktwxqfqKRjcnxkBGYHT+F
nhNUiUQuIJwFsxQuig5nCGiRmrckQsTwImdu99fLtcVoqi4xcexpUc74WTU4Ar+bTg9fKzE/BCxI
6aJMPn9KTw7f/9O/62DeF+EmyDe+0XbQ0Vfyxus4FigMs/rrMveGsiek5gLkcfsaCmSDVqli+m+W
o+J2i6Dp8nBleqfplFtBPDo3YlVuxGrx1jZf2ZYLb6t2uFmVKPSvkwaVeZV6qLzuEzaps7jpwZYu
sGdtRtIPjDC4QRq4cYJW/lKqnWwcEWj2yENtUmxtU12JyS4SO91QfkYsZC4Uzs25P+cbp1p6a8Er
CM3AiXTCvWBFnKe6woWm3xfd0SsCOWnWwM99dCcPK4Ue6NFm6MLpwKCXfntRNP+TY+peh8AfI8XW
WhITgg+0TX2It2/afj7aNZRNZLQHE7NkDGJxmfBI/Wz6jPvqyra+YE/sG9ZOK8GtkRtFWMsGhwEk
/5k9AUBDu9SvgvKYat4pRrbpcSuViSkcyhNYgTIB7xlOvMDQU6N1aaGY/zQznaIpLUtotqeWcWgw
IU7HL6uZlCeySR63iWoCeZf4ES5/lD2BlLdjv06jijne8dpQ5BqmYx557eTvJP0A5WvPcIKOe0F0
lUipV4jbsoffdCBu3uIRR6KyYyNBGvfBw2HbQQ2TbalEQb9UHI1QO8J5Q+2VbOnl88AB+xUtOtyx
e5tUmlVeuMGoYQFXjhrxa6MqYOPKk5Uq+T6dJVXVFGFTBoCrH6Vq03xKhsx9hZXaMu6SKpcRMa81
ahZ6nVwq1UuiNDn3nnmFWPPZ4NmPLH/ESCQh3xCqpcL4t/E3qqKAXHPZM4sWx4hKbJFDMMLjKXdl
OLNB3ItPGBrsbpwpXHhtbmTQRUT7OKnoFY4RIfd64O8wevml7EA3N+JmKXLdrQD0RvlpV8QItaK9
LRelTo4hWouzWIipemDKqTeaVCEJ1OhlaPQbkEum80dzUq4ZBzxKyI0FOTJlx/gwKiI3mJndNNXY
PsZUVcs3rbANrqUZ7fAsyTvrg6VB/0OPlurPbsFv9ZwVEWZBk1HHfQPbTIxAjhuWTHyV1VzLBEpi
LOfueIGaxWaOf4utUsqQyd9QW7dxTEye9z6ZwNm94l1PYEQSsztqkZ3YI6mJFyg7ha5L0NEOSsjo
sEUBvuxPIjxqLxbwprDoMMxGz7L1bTq55Q2QEuH0RI3ukXggvnc8UMSAMAEqBZBrh4WZGOOoKBRu
x9vM5bf2xn0aUtrq+jKLyc+ixiXyeh2ub+K8PO2pGz8fPDt2RKcNfFyiO1ZCivAga+dO7YLCU4mJ
huAdEtkidJ/oXqDlEEk2LvDPoutJXdvzeziOE+5Cf5CNHhYE/Fe/GIPmHdnrwqZQKHe66NUHOit7
81H1lObysu8fGFX25FPlWo/mWNUvJQK5JqpcRBQV/F1ZMqYaxNwkrD0jsiFSGnYnDOBcfofw9b+t
QIbgct+ojTcZzO/LtJ6OeFW7iPGhX6WxDuXeBrQ047ObAGVvl9DjJwPnt+uUPD0fjVfKLpy6gL/3
swkoa5FE4ADJQszqTPFgCBONK3bM6E2gEzeoE3wWX/luJnrzYn1r8Lv4xU0Fr2I2uFECZe66P7cb
bCeWh5R6BfE3FFHm+dB+kI5tR8pYq+u9baFeTrSITfnTmHDdAQ2z44P/AGRuHlm29LaqZFhFZU1l
lWQQouk8N8upUPZi52OPtsRQpJNsrM3ClFX5fs5IYRryuIPvC4uUmfMQnA0eV3aKUVoecHFWZMa8
7iZ1vPZAiZ8xttR7WEJJUsJszXfFOQuvCGWAvFfmPYHlEHOpC/OtewiP1zSC66Wj3AODLjtrDbbp
KKN/bb96RZeQw0xUI0JdWsmM48DGE65EJc7NIKHd5TyedajFwhSfQp5WypXEwOLFC/8uD1GJTcT8
1ldRB9l+M7HiZLkK3/bR/u1NTn3gvY/r6Hoe5B3jPT4T/l9n2Rj1HmuMjoevOJkFhX/lIc7rRXNX
DcGt3grokAagn/yAJ8lb8gKvDtucQtB1VZlDwkiNSAVX6RJm2rOP0z6C4agepuUKU101k4DPSOIS
sC8aYdYBHClyc9RetlqbTJWuR5c4gJvsiKi8/d4JN+1mpguc5Ah+eAMMK13LlvOd2CtIQZ6wwjh9
FtKVgZ7a1oIJVRRlwR1wumWiOEma2d1UMFhuv4g5kHpF/GZZd4MD+72pH7g5daCyLL9wBhnkyL+E
rO5ctDSbeyIPxL8np9mVN7guIQ5M3yZ0YrYIZ9ff4AGVFFX+aLLb1RWe8O2gvWLDeOMckU7dj8Iv
ALrjJZcah0vz3HG2ofNucHCglJgwouRsG5fIRwNReZoI13XcEY4uhkB+IkWKQlUjINPkc1rb57Kx
XHa9zxDgF//SZWQ6Pnzr7A3ahUj4mAq/7LG7W+WfB4+DIwGTIzFGIQ91sm4MuyIBOgPvCggDFeXd
XUrOhXrlekf1phnZQoCqnE50z3qEx391RuE0E837OIcsatyZ8Rrs5nLUcrWKJO6awr/YKNOwuP9t
nRqA5tU+OEdyrSvemAQ6XsCskiACzIla5q9KGu0yAwBvuMoyn9A4H0wAirD/jiKQzBrOf9tc7Chg
y1+x5HAsEyDF2+k7iAj0eOfkh+52oT9/2SkCrNpv4R6HjRX1WLTTqeKd0HjP4qTz1UhpnYOfL+4g
U/Qr5m6hF8Z5/kMl/jswjKsTEOiqtRVKHyKtu5Iax6IIdMPhjHhk9MWwR9P7oVoveYAgG+onMsmp
a0nBq5mCa2xwgCZGNRwoXo2L0wz3rgDaDrNyCQ0qBfBU6QSliJ9rqfaxgo3zY0xLsUYp0HPX2o4B
ppdQ+sinQN1hylB58cylV0wynYa+NEqdePqA+56oivTKSJdT5eGddYc2F50B0DkLmPjhwvrmlsA2
2RQm7GD0I1Hh5mjsfs1i6XWhUudMKnHormpxg2CU7Q0L5PS/Yt5EtBCpbXlnCAhZmqGh8gO6I8G/
Qwr2DtE453rL3pGSTovI18f4Zs8suRm+jOrE3BTcYzqpESef5s8OBtRAHMh50NcFpDdIb+OuFfTn
3aHkmwtWEdLsa+NVQx7rr+D773ctaxKTkfMOTgertNprTopE3ZqFDFZZ3I/W4KFPSC5lAVnf+Esp
aP6IflYA8cqnun5z/NTNMKUEABfIRL6xZV+9wYGFXcza/bNV+eU8fIAOUs9Boyy+4D5Bh/IV58d+
lTpEaT3RAzsZHnTOKWlmHngaybIL2kCKDuSE8wM/B4r6P0GF/BSy9jGm0BSgdV/7svSWJMFe+vL8
3lQAV25jqZ50J8mRKcweHU1hBFX9f0iNCYVZykldN0FemcinY/KNTQ1SFV9Zt1FVCYTlcepsGPyb
LJKbQ2UVjdYswCN5emXzXqXZ+n0QfmZtkFFHT6ARxwRADIqwLika9ZHbPoxh0H+TI4SKoGBZi9Y1
F49jL9IVhpZ5TW6VzAgUHEt153iM9Wan2K1xCFdjL4JHTOxp5pX+jfXzXVmDmbb7CR6EqekYztGm
HUFAl92AdDipcpDzUCIAr6Mw8q+mp89mvfCdboBAzXJjHrpxsElpO2JM5tZM7BptdwhDGMN/3wdu
9MbOPo1W4EJXU8zGRgXjoyAXvIfcl7rfO4ZW5HCCoUx4D8rx2Bt7HoRpTUd0IS+NP8fqeS/a3lnS
Nh4AfRMFCC+1ypKQNSdIF6wp6mceW997HAx/twfpXDPJHENqnN+4vII8TxX6lz3nOOS489j8myVN
RhB4PcAXBE2Ezft+X2il4CSTVUOTDiNzqngoEOX0t9hxeWzKpvDAZv1k0fxylsGzQdnW5wlhTWBI
ZGJZJ679m+0F5Lj5zTppTw2vxJliQSeRxiEZYf9ht5eVfSoGbVgqFCtiDnndM2wNLdOFK3CaZnLY
4ZMkaY73aSwU0ziYbmxD8+Lmc54R5/iJtNDYNWENKnuw6uZXrZm4Q8UMc/7f4qfLSfoErm2hMLaQ
OoZHDyaYMtkwfb1qd2WrDYwcSydq6XOD2x1BFApGAaG5AtHU6s54a47AM5yys0SW/FpcOgyjPV+I
2ojVyz1dXNeQvgr42TvzCZzFlce+IVyl3JgWDezOAQasCKFOM6Kv/gJzsOmJdZqMhDJLsM1LzNiq
0ZNB4Gi6kHw86VPx2KCtVqdc39TyOQ+9xvhjKHNwclak42yfnsn5zwgxxcLxlvSCfr5CzLwN2tsi
a3YjVIHCCQqzDkeG0me6p0T4vtmgJ6gjPWFcrknnM8LqOckVqrhyUhmpQxNstRRKSaXiG1EsdTaq
1QW9266+5sAHIy1qy+7e7nb0kbCJ/150ireys9HOGZBRLOiV+roVgn2UWyEDUjpWBoCFseCpix2M
faW/GDQQH1ufmot9UxAdMGpb/xja3zrG5MAcDPqv/P9QUOukkK6dWeetrtxAiux9c7JfHxcf5pZW
LPIKkb4qJqJ/WqnAs2K27dPVjyHD5S++ceEuf4wbF4uKw8nzeZhVmOJBdYQ/mIPaYtVXcaYw06Od
wb18Vh5+9pjTFjRF96NrV8y3lvTi+S1y8okVLy2K+fi387D5Tk0neIYJ1gwxGoeGKDm0TR4WuiPK
YwVFPdjdUh/yHDUhMJ9Plq2ZxtRUO0dVNfYDKuX9aay19LT03OnOc5bycDABkRogZytERK/BcyMF
OI4B4uW+70zp10hmx77OhoTiMqv23ocs4xG1kfWTCHyq3efKsxmNNIxZ7uV8uA5AW2tGa2WLRDCX
4oOUvdpmAbN+9FWBZAdwwRDXK3d43RmSFLVqs9YxU1Mva+tzlIcxtfHHjgYtyM6CcvtjC7Hnskci
ZdC75kxuhOS1eNkYx8zvF+EourllNyzHbU359Oxz+Pqzor8D87qZlvv3SMq3QBuQgglX97Pd7JsJ
HArHooljg4zwfBvNQDQS44RwlEd3X9IR/ZqzIp3YgiHfIZw8x0uXEK1TclwgMMM4EZAfp5bEpXGs
7W1lqkKtOXev2Z9H76i5K0V386OwH+V04PDPJTWE2c4Cns1rKsSfiaqKVE0AWvKYR6RxAXyATh0U
MyHNJVvytuGeCVrFoCf6z3segSbSg+Mnru3xz6OpnrCVXLMM8KKnFh95fumsoXWrxDR3W5FfyNI1
bAxUl1D/mFFuhKuNgKUdTu+swu2nfbiZkHhUc6E3jwKjVar2K2uoGnmiXBasrWTH36yUyrU14OT1
Zpn0FBqt/uswCPtfFG1bdieqlJ9LJ8Ae9jPTED8LvlAsBxR1J9IMnbeqGL8m1+LCZdBBvx9mYaoF
+niNR9SeIzRp4plGe8Jw1w97Im2Rb2s6jlY6K1A83kYIgn5yuAVtk+k7JKJkQqSoSAUVukoLfeeW
Li5PHwZnNJzQ4tC+UiNO+reqIwI4qt9ujxJSI86+FUsiJVMfbmX+CgQQ2IxssBuUveV+g2TXxlA2
AYTs72e+6Je/DTYRFmZW22vTc0fFcOtg9mwihzbaMnpeIMSlnSnyFING3imti+zF41p+eGNyXhpu
Po2hD+B1IsH/zVrwW/UBzqgqAyVQgPGLDvVTcXu3ADQS0X+FVIgdSeEI0t23FFqEk7hqBoNnxgeo
GkQtMBMXTq0R0AGRnr+FOwymJot6jsQ29+OehgzLPfCBKml8XScVQRYKvOxzyIJ94FyVHLfeL5Ih
L/lUqvOBZBpwoxRgoaB6UYBqyZkuZjQZl54HgTt6MufeFOlJZWbiF0wkmjyKLngD60awmduxRWai
l/9bGEOdgh+jXU0TaBWUzFWUkShoAQWwxtzo+arU4QuCQiTCi25xg6oyi0JUkP7DSBNLgvzGHFxz
ZuA6VdyzgbQQoUJJDtFmXwafxWR5viLXsjcVFkquYshcLrkIr2MTZwstTrl4s8yHeBvZ+aQ2JqNa
vo8vrejQ4mG3OJxt8BlGqwAN/ShiAe0tCRrvuJ2Kuqbtsi4XAQMOTrCwmP5tUrUThuvs9oVLXLbj
V52vtzKZprJxa3+Br46om2COH3jHhbVmbC/9u3LGua41CDbDfoHYHv2LPFVhv0Z/ecLAW+zvOFkH
gXOgS/bDw4BPfiJlXUP4sPvw9j5pg4xbSqJaviwFw1aYCM6kOGz/VBmZemER/HVlR/gC/M8go4jb
mgAmq7sAc3x46hCr6MeSELUpR+ZX08cB0NyNlBmGkTDQRwu6+OlTkAtLTS6VZS1nbC74ym2bhA69
Bu2I8efBMZKDzfK98/YnL0OwbvT35j/XFnq/aqCVbr3fqbEryXhUiwIII/Xmz2TJzfcakQtGb9Ay
PZhwi3+KyBt9PICrdZPsa8V3p4OGGGoCseC6i+HLqJAb1/v9Gldb2C7GU7mdBPCehBrk6aBLbOX1
irgpTab7BiVpcBO3pEDE2i6TWQzvjZukiBHwqcvlg+k3QSGRoPC0wDXj6RrJVNn4UBjeNCQGVu8j
jI0ofgYFjdrk3KS/SxoPlmJQ5639RFwV1N8SmX3LvpD6zeLijeOXXouuERpv1QDUapQQZH1so+Bw
XVG2woKIgC7r0k8O6sYgbhSUc/Bbj+OdetCGqtkRAqxnyUnvzStjXFtFb1NPacShzEv4dykP/jdr
KjcWnb7fld/ADA69juwPWu7ptwJujlQxqZKCCHv7Iz4JKGR7E1xKs5SyEwR3SaNKnt7mo8BYLtOC
stK5y7LN8QfvKlNg+ecKjHZjw7vIhX5k0SF6LpyJ/tFTDuBxL0+6DBtnh+che749U3KxS40HsxUa
QEWEhxAMFRnvZu+OrpQR/6/iYvlK2lVKTrEedKEYv2uSGu/3E/tdiLS6NEGq9EO48CItcTWj1VT2
v9obq4MdF1b1oe36KveowsCmJi++7SH4162hIXiNSCIJLH7PBec1tywlax3tByRbWy3efCF4Fi6d
aH8/9tKCYSnM/xEDLVx8T0T7RDRYaeZft0xCEr7YZXZxLOarohvYPItV4zldrEFchAwIlQTw8fD7
OwITdrPqSK7DSRQxwlpEeciFj52YzbgXUNLOANdVLmzJOInOmBVrgLcUUhbiSs2WcIGuwMjW2MIu
jZA5amJ/F8jI2XZLgeKnK1edbIQ9Qkfi73EF3GESeY1pR5vbDBslO7gF/n0sw22Y4KpRpRVxjmgh
5xGpg7UfP6oThBk/vEnuxrQGNiOFXCblzk+RTRg7TAIVD4gBVFNvXhY++MbDrzWfVL6hNtHVBD8h
MQGxog8mNoprhyiDccnFu360+2RaNsrscs9DylgcSsXgeQasRq1/8Er+iKoYpRtjBVk8gtbcDCNS
Cj0mTNry8yjL1zclhAcHMaWqer/1RQtf9d2MCB9sT2aYPqu2LGSnYtiigi4GJqzgdU6Z6cWpx6aj
V6SePBf3q5LEHIt1dJBcmgKK5az6mQroQvrfKMG4giUte6CdZR8qzIomynh57XsyfxsYyI1d+o9T
0d7x7+PzwSivMlKFBLMrL86a7kqT8MRH5CAD6NP7UOBtyHaeMVs5CM06jlWnUH/nJtbAvu1MOhIf
N/GVqyCDg7xIQ+QT1bOvwGutMt+DGsXZGNRdbe4kHuo1iEdLrlGCNgMxQOlg+vF7BklwWJeEW0MZ
01xwAvPnTrM+4DsM+FKZtTqKQdTCh9j9L3kp8ukZ0nj8SfePq+Bi0Bc8prSStEVfw35sfgPbKihT
Xm6ZKuYJOBG0oQRsaZUafea6g3XYvfCz44JDnVLFL5NNX4OSVncGiaAkgDG81PuprD0JaSZqOoUK
/aeK/j1V6S9b+TYqsNXd8Fk6+mN2nKhwnp3Hyg4MrcWj8DcCv7hFLQdqISYnqIgY/jZgaITewDtV
k2VaWDDS3JkFI/PPOIyZN6e9oeZr1KyW1oKZ4DAcxAk4TJcYroLL8LGBUpPryqFoUQ+4or9povCf
L5umRnNgHiBpaq7ePmiuS6u1yfftYLbnvjTf2DaGsIh8aUCN8Ia95PhxFktGw9QQFN9DJ7JsHlco
yBpXmBQaO/cIX3Hi/ZCBmpsABFKSErHHn8dhUUzJ+9u1Bepd/fVh4EksqQRNjfYwKPAgQ6VndaGO
KWFGGzGYWXSDqZ9x1AEJvs4fH4trXU0J1A19BItcUr9CgEjxUhzwKvkMI34JFbO77rQU4RkBGO/Q
JT6Xf+a9QQAhM32Th5nWBi5xIh+sU2bngkBLNSAuhg6BQ9/3nLSWKPi32n3fHGAO7awqcUZjY2Lj
szlexFUiFzP9JsX/n8zz/UwmqK45rZ8fWIQYoBbmJnNeB/mH9B1FPN3f0Zfe65Z6WkcmtOpVW/TY
YmbDrI1ZewdF0+bZMFyhw+OAhIAgQkr0ZPs9WxvkvD97CoktWjXIdeXdPKHr/4+2FRZ1OVXWw0cu
7ucHfCuEVO21qakomtkf9ftOgc9r/Z1xqyhH8VuMg/XGU3OS1cqxcpF9ISXOl5qMLPPQy3cPiL31
vuePq4pMhdenV5zAJYwFHyKZM7+WZIb2eRXavxoLB/ZO8K9yRxOI7y7t4jGOXkGWjhM1Uj5vJwUp
2XcFeSV6TyNmcEFB/NOaBK+1WbUATCmjI+GPv5hITcHm5gTAThDb8SJFNy8ETgTePfQSe347tmRf
1SiD75RglI+nXw3B2f59zHcXIehXoaNsXlbDGatA4gZm9SukXpv0mwPsq6qc/zuP8MFCnhLKaH3E
K9268G+sMY8OawJweLcdRCiSyjgy+GKeSjgkbGF6QaVHIwmX3OHu1YhK6jICyH+oEpfc42Taj+ko
Hc7ldWvLn5JnsgTmc1yD694VNItJ5DXja5w1RPzuqeJOfZ6IV99sa39Rb/usTfqkGvMWsF5xmFiV
/044qCP9oAWVirLPiSYd/N9/4ldSCwKK2LNK1oWpsk3jcFveTTfQcg81b0qqdBqxjOkloHkVUv6k
VufB4T8Ix2uxkNY6bBmrEpRUh6vhXt3UANpuIcplCs/93df+mqliB6ukpIlPpXTwD2EZormyJGvl
S/Yt5NpcSsi64pEIxZ0CfoA65i7FAeYXVf13KcBFt73tY8SYw+jk2/XtOWQ8UfzlTa3ZRFummwaa
SKKpG79fDmBSvQ7kmeRfoXHTj62X3GrMi7amxRf+7Q1filZOwLijPFXpGG0ykjBNkck/TAoxVA93
IMiun6xdiG4Md+P0u6KRuGcg8GKcdialG35eSahxX8BFQg9zzkc5TrKFfl7yBsDrXBhDK7mPxiLV
6UrMp3jal+SLaKteM+MjspkoD2+m3ilBzGWQznRwga3xUJM7bSiz2kF0+pQBkwhTSjJX36CwvHQk
HPTAzwBilzYrx0n5EvmoStdmSXN/SsHNZH86Rqd6fMAemjFSD3R+lh1F8SHXFVhF5h/7rMOak45X
EgPmIB4VwF1uJTRf1TN/8io1BCWHauqMK+MIb2gk+bQW+QrGNVZXj0IT6Jci73dUYfBTBsh2Ggae
uH1m3ybfa4pzhjZEvwAHr+pt4oXSE+4iRFts5fDSZLZKLb6pdCRDDXfEOGRIHBUnKFUPgJ2KJ03Z
EWzZzp8VA83FaSk/ffIFinhIRIIIzcNwdZI2HgbFsCczKVgm1joJWtFDOZ1D33jjpxFC8NSQV7T+
TWvVho60DTfetvf+2djYwFJUze3sc1ReI3/GdSMWn3JWnuXPTJ9/cX9UbkZQOCEHZcPvpq1dDRCC
yTYBVBpofkaFbn3jyAndsWQo3aMDgWVhE1lSQVK828RLKXsBHEHIAkTSQ1D6TZ3ANbkmok0fzuSH
JG57/vb+9bRr/D2CugVH2HXq4JZvhjze02RI0GFhQh6AtH3rDLmt6G7B7VuZo5YnRhOvhG0HFGKx
gOoThlhsQPbJmL+wPlPwLc69/n9YyXJDKq99XoFxWT574aE+9ymma3/DOxfAgboskTLEy3zZJSN/
5fXFXO9FITnTfxYgyAUHO/b2zdss3O1w+9s/KlNDhNw/oEw9WDhSO4DiEV8K4ezevRA0750+siMz
N1LAXIPpbUn/OIcsGrBiIwBWTXJPFYyIyn/LREQPaO+TmAcW3UcMmifC/GSe8YLLJUT4GpcHfW2z
RU+NuL+cT7xaLXEG5lhf5onNat4rUJc0F9lxoChzcj2AiDNAA7/E8ubrWmVjnXoMIKzv2krlaNyc
1URO38XpL9jRc6Fdi5d85xHWBge8imV6QfNNURDIAdFVgc99+Rnqf1sw1aVGacWZaSFIirHodJ5C
ZDY0VpcQtDd78+e2QmJ4u3kioaUjB/Pxn4MI0119Qj+ebtw3+ZJjVGVnV26Zu8aq3BQoNfy+IsXT
QO4EVOI+ldiktWK89W5yx0nKA8BkCJSc3suY9ehECaAQlCDM1zU3fBehk8OZq9tXu16GNuTMnM16
JobJkk7y36h7mFmbkiOZUhUrjmZp2rCtiyGDJGf5afFl3UyfPJPRq0j9e/1kDwdbPHfru8eQlJ12
/sCuTHZd5nJ0NeOWvL+Mg8oq5NxcFNxDwe8GHtgQnUUt11dKctuqKSWloPZMcOpfv9jAUs4U56+c
OzAGtzoseS4VutWJO70nQAxs5MrycZAlCgJ0FwwmezFCvM5FMYRnqzUzI83q8aeGEyIWsOfoURnt
k4uupn49dcLiULwIgEdkxAwbtIR3an3haUvPFld+/8UawFjX0K6KAbHM0UqyJayYYn+lK7RL0BZH
sL6swloFYovg4B94Eq4z+GKPzTmNTyvEtg3mOXnyLDfHreMzL4cvFWUiJbZzbyEOD0RowL5J6dqp
6k+T3YHPKdJxssAd32bna4OX6V9hG04ehM2cb2wWMc2oYJ1F4zsae7/PFbNPEsJxdojInuP1ALzh
zfO6N13+IvxMigqSpzJ/IoN2gwMuT+tTOX+wmZVtyZAkKi0t6FSDeJeAfYlaJX1nLrMWt6p5s1Ym
EgOsid1RP6xysLR6YlTAE/fEiBXYsctbUa4SzzhNqvkLst5I7TByDr2zCxpF3w9A1rd8eZtRToDL
A8IfQJdcUal+b2X41MVmIUlaecsfHJJJcH0pE4/wWZg2GtugdG/g76s1yIWR9TjseIzANAGaB8oo
OkhwyKDl9huGa3hGCMQkBVqb1iaeMamHLesY3bGw6cWZQCmtxcI9PDvKz21K3IJKmVLUNNdYH1px
/AtlOMGLfRLytkWexXUQMTSZL3ycVu21boPSQBxOk4w/AMjE8y5xyrQm0GPJ3D3b5uXUH32UAdbA
ZIETP8UE3DY7LkehbCG0+xdWMffR4d0TOhOFu4komnpLdzih3mRXZt3r76fgoD40Uv4H7R5uVQWd
A62TCXEYwJwyb21Wk+otAUrd2CdX1UmiIJYLXn+msAVM8wDGuJs9fCRonmwmxtK4LLDHgXHzAvmv
nzySILfAJclIvK48mK8kc5smC4N9CP1RSABMFeN7cDCTYrX00aidUKzbin4TABkcaSjiQ9p1QRJo
C7QChl/dC8oskcCmigoxcucJL+o8oqkfcko+1idcwJ6p263uDj2/w5aYpW0OyfG6QqARjCxbZ2hk
cOIV/Rphdx/4jjc5eVlcGImTI2MaR4UpZINk/qK92jtdpxGZrinEGKz3DNg18e/xMzsmFiCo1uVM
ZKc9ztpFK7VxfABrNhgjKWF2PMXYbrorhDuKJctK1d6BuLc+61j0fAQVEHpkUdvi9EH5bukQ07kH
O1kh2QmhCrjWDvl5Xi5rTgNY5wQX/dA41tHBqMAZ3ZhD2ZtPwoRmSfMdQqk2jH7cW97v4E2M5vGd
Kl9sqFly/JfKV5/zZ0YsS+dp3ZxvB3yOpGbt056FCG358mltzpvqkwVXip5PoaNksAY5sZ5hDd5y
v4H1rpX1bXSIGlfEM9SUSv1klfqUq8PBaWxstt/2H1CrD7LIEBpBaVl2EFTjLIH3p7UOP4CuXYms
aXb7bdPwBVqQV6LiLAjSCbhipnNT3dov8zUTEzxgbmJxXQ1hx3UqmvixGBsJPiDV1YJ0nPxiXRmH
QsQGgWyB5D+MJzWnzypagf3gJTKz8PFM/fv7Bb9NvEC/hcR0zvPgF5dP1GnffKpLufydh1LkXWdM
pdlAU7WqAASJOdXXGF8zzBMsIt+dCb8pipFEdXVD3cLzbFpt5WZsUBtqIeLiKO5Ulp6+QYt8vFx+
B/E9yqhWdnFPGjQKwsS8SeJ5NufrwGFFX78VQcmShPI6jN8yZt4dEyB9c9VvlmW0csKhN3z1tfQL
58t0Hw4M868NlyuY01K6IIjLm0wlavryrPDVFRvWW3iw59af5+39x6ze+QGRL1HoIrud/G3XNz8M
yuW0OoVLo4SLTuOgjcJUO76LmQ0wfOoUuCwr31ep1N13pC5dTCsf8ULLJbEsnLrjodGF5HcuR1bT
AVMZt73BrEy0tv1/q1InPqBNckRW7vuZT+Wu0uOPADx32hQTwMqFS3sxo44TNTEcxWPOlb4f5lJN
Sj620jMzPGzcK3VfNI/LMWxhjYvA8Mo8UQCfmx5gr0uT6SgIl01yL70HnZs35Ok8j0SkOHbiMSpg
bM5vlaJsly5bT6fZBQx62jVD9k1XPb1yqXXerIM8+jW3SrTKTRSjfKWHAxZk8WM+ALYNkBU93zeb
DDam/ffqAqZQqIz8R6L862TBIuMMPM5ApHTSGDDbCoI/aI+/40A8P2sS4AlaXG4WTStfASQ5W2/+
WJCgWBG5kdXriKbW8XWP4tbEPFbWUnASAlNPzctXElrj761B4VoA3fhpnrCeP8pZCDXX51aHTGD6
X4q8KjLb0RqEQ+NUakc17JIjuC0cv7YLChOGsxTUQOHGxzAVy4M4cAiUVraeg4JRpYyJr7m2DEhT
c2PUit+M+zWzfs0SMbdOKmhEmZaW5ZLGqEVYC+dLU5joev7og4H62kz8kYj+6sb5OjrNfS8UOdY7
xvKjrn+c7PL8GxBuDlZjy4etrNiUgSRb0cI/tRM/sFY32gFWhqEF0yYjAOVc5iCx0DSRrRBNwysL
HEa4kfyd0QcqBf2uLi4OHuhYU0iLJ0AmzNH1lsSZWJYW4EMZ/0AiSYtX2Jn9xgUZkBTcEfqyFkwo
C8MGjsMQhC8nnRi6jrC+hpjNEEm7OOisf4wUT5dbeqiZ5vTNivl6php9jNiWy7us/pqUJQnWBPUM
CmF5Anwuv076JLjaEinfUtEc/JR99NrC4FjyDA+vEKH1NFvdIDvLoqUJO73qXzFQrdA0L8+G9YRl
wm68Do5YYm3pe+vv8hBLAmdUlRedzM8T4UwtIBd8NYT4zvK3H2fHZBO6AdOOTR7KsM0brkum9Q7J
4w8RUh7Tu7GinRhd7HMs7wxfw7nXJ5ahuu5fd83ZGZq8jKUJQJupONjQ1aueBLIM4AZvb0+oM5gd
zfRjerB/b2NbT3LfIWG+G06hySADTiy9ReV7r9BS2iP/5/pgMGaFYrKgqnLJf+6KeG7FbnVGZKAl
Vk8VMX5lbBsqronOQ90o+jGUZu10vBrtRyKxj/vND0fNM+C/GmHa9QxvEtMln4kfqvcCtu+Diz+u
zvW9/0jaEhnCj32zJywOqTTatbIPV0CeA+CSCD1w1jCmybttzhJQX0FPkTG7czClIJGP+jnBKbsl
f98HYzflHKwTw2sCEnNLfg8/v6ndISV8RUhNvqzV+f9LIzkr+KjOOHISGAaSxTQNwG+ss9z3hQQS
N+d/D4ebEhqxBCeojCSKm01cF1x72NCzBNREbJjOcyRaRYYRyO0Krqg7NfsqmsquJyWIXjZZ+sUM
BppZdxsw4sICoHDpXXLqwL0zQzceLi4sdLfOSRMFU4Us4rQn7HZlVvTKm2doAauVRMQk16MVvw/8
eBzdx6DqWP87mVfQbtjVTEliYkneUi/SDrqsLpnlgKT02R8N7fX12SQi55K1e6YoLsLsr4VfQeUf
5r1/VadJOh2Rev0AJKDyjg02hqd+4sGnkrNC6wzG87BPmLG/fqj1oI5Ow6cV7AWmKBnX+EVMpUuU
/E/8OTKjzR657k9+/ZZnTfA8h3yA6zu+ixD5sBor2UoENiaRqxcin7JV2dl9bZwTCgiLdgOuwNYC
dFoDLGldMpNNbdUPEeQkdSGp28A8ntlM6zJUxeKbyoIXkwoFMBefw1dlMGCvVM5GjNQAx4TZo1WC
FhjDDDzPTfKY1LOb8fvkxvp79nGzbvjI+r7mb6Oko6Cf2dwPMcGOEWVnwcUWacnX9UufUkA80I5z
iYQ/QqzLOwpUjJ8yG3SiAU8DT34NKeGfAMqRfnarsiCkPxF41x3nqKXaqmimI+6ZblsOwZkIr2tZ
UO/2DrmxWlqdR/HpRh1O9rW3wKZ7qWeSe8LbUgPvYiQ00mnGMuKdZYH631OfTh85kUSdAU7eH+k6
wDNXHWylHDXEBt5kWjnOrMUQxgZtougidbvvOqrIXPXRaMZ9q8ysh6QCnn6qCc9dXZUV7g1rwDqb
pA6iYQ5PS/3Obh9hKsHfO4bkQasV1e043gNNdulDGVraH8xxc8D8wtSlYXTUjOkVIg0vH6Gj9Q2r
Ms3VTX2d6Y7WP+cFt9t+nVG9aLdCeFm9gdbwT9MKWSTicwk+kCo2oOw+G+AitbQOyLT0xOfG2s+w
Wble/64IYkDN9zzjL4k0LBHFqLDMmwvcxyMvHFENcyqSoIaRIbpFWp6Ese6V4WrAXN0ObJA1Gu4P
qI05suUBSLtkHpBuXrL6W2F66QKewigdrix+H+Y9DFT7DJd8TZzoNkC8OjlbK5ltzLEomJlFu9Mz
2qy83irqbiTcKgEXG4+lslEUknmxaxfS1DC2ppLx54oXwgThOs2ll0jdkPEAP9ESXX5mRZOiypvv
9mIvNvwqPY+7OF2rxAo9JAwjAfa7OZqKKYDU8dsugeY3wfLtplSxVQtMKcgIxu61slGWEm2TtV1i
PttQ614HSCwxqXvLkMQvk+7MS7pMOtgnAyL6GTJvT1tHNrhhwsNp1CnZUyORu/J5/JLaAZuCI1qD
j8ypYpbW8izf6pNVmNd8ce8Tc2qDYLmhczF8qO8pUUOjqvlDlNzZHX2se3fnAPVdb3bs4hh0qe1a
NBHNExws8VghOEgbSF+35NGphwreZbf0yAlgPILdMClxRUyz5Shy6BTqhq97+k95AUjeDJHqVnfI
fQcLRBqZaIrZg9jkeVa84jDI6SKtdEV4yldKMgAhKXIGUVDmnCzlp0S1yOnfpoCRYZmHM+PhqAeR
BKH3utL900xaRkGcVTVnTpuclcY+crBDnnbXQR+NC8VbgGUlIWulS0cziXRKjaqNSJC1MDBvzsAD
2U8QxkmohECJbn0wgPpsUybScu+GDi1YulaTZkj0rJRNEosWui4lHCKZyhy6t1v2Z7LdXIiolveE
EJDbbeNjm8YmUm9I5r/3LwtRbOOnOfsEPlcKwFWv6+PzvEQG8nBWbrlhhER29/sdr5KuGmaFiPBp
IPQARgZPbyJ7EG5HBa6MeqlpcNBlli6JaYiZpDHHE+j4YBPwCpjvRUgirL7msLpZRdpXZjd+1jFH
GZmQznFlXwSWFfcQbUuElruAE02yi0Uk8vOTHsdmXx+GlYrvH/B9twok/isUBJXiRxmxFcE9d0r5
dbL7/jX2hk4b+ooYE3TRoqKEJZPC2YQ1W7o4OH+zejhqnIo+hGmm9IxpYZAJJRWiiuHCKWA4MHWc
KeOrA7GwePibLzzGZRorzcpXZWVkSLmFchbY8IPcIHGgFPehh8D3uh2chdAY+fFb++Tnbcfh95Aq
E9tAIqZax2Ue8TPp2AYBNDTm1E7sninMt3GIJoOFJlZ/oGuKAI4a5wW5vJdhPCeip5RV9Zudg7H6
GBA9fDpmZyWgCFiQDM7cescUna1d6MuMjPEQO0zXeG6OmaRgBT0tdeIKUQ9YDsYGjaEjMZ45Ugd6
A3LyDILBc63lZrWpf7JFFQbuEMM15kDvXNQl2+GaK8TDuRnUVI8EJxK9Gqw4EzjGeooDKgWGzk5X
Ig6J+fc33KB/p6MqTWleqtSYX+GxG68Ei7YyExgiYYdUFs6fcBBwS92m1AlFuQBsCjh3zVoz94h0
7j3n6u/yELtVnDcicGkmb97m+Jq6sPBUCUHxy7O1v3iOt0huhVI/9Scxm2j1SgYrLgmaCgQ3d7BM
tjGTrb+TiqUAtxvbns7fdMjjzATbejs/y7JP1P+uuHiie4z6Yhfhn1Fmd1YlXFKJ6j63SBCoAQXh
dB0k9bvJw0dRhQkw4uC/dsmEI67kDdS3lEC9ozggSkkD5WsTZUKr8kg0zkX8vnwsCodqRndP0dJ9
gXLDz8vdiPJBCx1pobApS9V9nw+KZl5apXUAgYOSg1Hbun0V6iLa4xOI5bgnHaYS1g+9bZL9Z+3P
u6k1LkrxrVv9iFKlUt66LwxNaQJ3Ca5eXRH45r2kmGDKCQyERWWVNiwjbcuMYZTucfO5daQ5mfhF
c2ZkZ3pDFh48YrRyb233QQGm7QeC+RFcKjnyzuNqWu2g/fspmufxtcahgEDPy/hwWPFqXLUtcPf5
fZoHgtvoicME8hadqLjOfjMk8ah0xUevKKfyGGp2c+VJ7zLbGWbE5kzO1G/B/wNwmYNgC0d3SuiA
UCvDarzXFhif2ska32yjWmlL5blRA9FPJqgc7Ymvhb5CoxRR0Ey5ZzjomNqBsEQWW1L+mSg8/dfU
iSLZybcwve0thBdtWiDSGHtvqh1Z9hWHIz7Cs07UHjsmaRSLmXaj7MbIT4xE0teJQlTdLjdDGjR5
WzxmiG/+WOqOuVo1zT34F12Y86W8qlRQQgushvTmukTJ4GpLebnH3dWqDlbLipvZAGemSprsLOx/
kCSmeJmWrlAy8StsG79VRW+AtfGceQ80wSahjNw5Udb+jLQJlPu5wBh7OtSj5XrLrKQhTPBRPIZJ
/nZCyl60Wt78/ow393/+65g4t/+dzdecng4N+0wMkDjtkSo5tjbPokSdj7U2RpQoEkSPnANvA7hc
W5oPaAk7k1pt265jwjJhwDEAP9h290eVwSgmo8SagNKsv3YUciS38NQMRJ9UyKKOxa6O6v6xBT3N
FJs7X5YrrQPAp3nvQdxiPlyqgHAekLjsIfZcIWAdcocbOQEE8D1QhWg5Bw+Ue/KJ+OCr09va1AGu
7Q4+xz2WpxBLTM1R8TUYdCFkUCH8cOhi9OKQl+jHI3GwPMLcSK3D2Gf3NrXjGG+BtoTeAl0hcWBC
Yi77hTdUg5nnNHe2pQx0wU2nb0gt5K7HiZYWHeylykmLNIatlvsySEp4UmwEVjbMA2Zskjp6gOfp
zXV53tnSD5K7HaMxcXxfgxDSzLQ6l9qvfUwNeqoswt5Sf9R4W6aCDOECbKhGkf3Cowa4+bbuqDkY
oCGrTZHEcmN4J6dotF+a4HjNC3T8yUlhAvcj9rYv0RW3wiBECRuIq5Dpyc5vkaLyi67GQgI62+iz
NBszCoV6DULIoPGrpK1vxPupxzeBrAR2v+lt76qJdzUb7deICC+U3cfNxiYkfPNmKc9zRKKvvPMN
5dMaLVq6c1K7Kv9DSG9/nNr4ZSAOXldRTv8c9uCEivEQkByyA8p/Yx725rR9ntciM7TGRp70ZYYr
w29b4ZGh4vBHWL1/M6xgRkFJ4B0AbXbqocH2QRUYmwKS1PIU7EL8MVC/FwVBxaqfWfNPJicrgnri
QXkF3j7WasPrLiI6nEqzBg/BOliC06z3BlmAGGLIgq3U0E7CKBCJu7GDEZtUiUEtskfTRRGNcrdI
lU42ZvFHuWmwlutK0Z6ZBubnrfdiZFYb7X4bJIPQ/zOShH4bXpMHSJxcXGzOSBk7pCY97BHlkCMk
oF6orQPQGV9mz0L31+REDbgE95A0waZeG/aHJxzaPvKI55sn4oOmC/UokJe0PK5NLP/N7tmerA0A
Oyvi7HRoVHwZWNgznpMw6hapekRLKoylcd3PykNac3QCQ3dTO/T6i7wKGmJQQIEobTAyISUqF/OH
Aa9w1kv+k37FGxozcK/itdIsDS4MC42rYm1nx8uTKwmqoPl65+4LW3FJApBsDxJGZ8QssoX/1oTQ
lwCB3U8iBMLjJ+oqoTEGTQRdF8JNLbpuoJjldxht8j82mr/CjfmXmVDV/ZEni3rfMdmoOnett6l1
qfxt/2ne3KQ5O7Is5jp68DeRRZa/plbla+2MytQ/q4KPVHLshRgQ+OhhEcTWvl2BpLwYODpyJ/4C
TZTlyoqM8Oq5zTM0cgCMQtk0S7NrQ8Kucnea3FKDsd36DROvms7O2GFVEHM1Mgt6s2OLnsVLz1gp
lnpA1oPQGMoRCjEPFeoXDyohMMXAXspZT/awFfz6lc4GfwKLNVQLarxIMzWd6b4iDksqU0nvvwfN
OSWr6uLtxPCtkG48xYy1n24m2laNHh8qSKyhcBDTKx+Ulmv/kMCCu/KO+sjAvcWmN5ep/O/eO7g5
DnE/RwrCMCtXY9nMxfmrObVg6VYG6w//AV6mSQLdTYrGrMWAQIUZgnDQuivewfJPAxZIJdvfO9kt
3Lja8qQTl1Vvd1L1Q+rXUPIqWU5Cy8oncs8qMQGqynMR1OSuIoWc1wS0Y1XsaJ16FmJSKqLvrdUH
rX1e+wCjLqtodGDOB8nh5zVNDhNBHTOVrZ+LV08Ji3v0Yo8jD0RBM40srsOXJbbdjRSe0Nq+Syp+
uL8UzrnMxBbPxK1smcgl7Qa9uNTU84lOxLG02t2sCojVjApl+Jd+9DEsK6cT3t5VkjamJNtTuEmB
aIU9OGtiCIIu3WCLGxlafYQpLeQccsIlD33hbL/SWxdabpL3ObVTsCTsh/Waoso8a8hyfTmP3Nvx
QP4FLBsxuD/+gwMrmDmeQ4Q1T28u39ZbW4pb3UXyx6b1Q2JBBBBHkkISMIk5g1Jkq7Zky+uhrABt
695QJraXITZa7f6/WKjteXtQsKpG9qy+fJFKlzvG0LuHCO+xzbmYkfwh3mwfYlX4wSNKXP1M5AAa
W8ZVcrowtar9IQx7C9Clj54GV7PO7vCvi32t+HFqxndBEEcAo1Q/oxzWFlUGySPqirNhCn5fmeLv
E+ChpysxYdR2ICfhgJqG6efDN/kS+EO7itPPvhbeyiO+FX0JC4YYa9gSDIiGn+ux2oBV15F3cDwa
zGp19nVb/CUPvODSImpCTYexMfzqarrmdo50hrivQ7na3R/+p9Uv4EzcOp0t53+EvYBwJkVDGI2a
altKAevGLk+oUqUqdyZhTmIiDcfI7Q1YXx5BgGLAEi0sPoL20e10VSlE2Z6+RoAs1ZanSfHLg3YE
q3bfdQbjULk1yjsxJbdT1ocl7VWSuPeG7wMc7sQf04J58WNCuBj/Kk+qnV6A47WK8vAe5xBHb1X+
QQPakZUT7yMjN9+EP4tFeZwmozAA1t0D214Hjdb6+mi2uYbd6bCTR7JnA1jEsumNhIZn3FCTXliV
Xtks3cQWPsI5bvmb5WmiTPttQpuWNO7xaLVDtnXFPBi80gtpbujiNzqeWhOdtGcWxLnNhociqwyK
Pzu1/DNgHdiApPciALUHHd/3kIq3sWqaWjG8r+/t0B+8r1CaeBVOZcGK2TDQ5I3/1MlCpbkCmrVL
ak5lIzj/UFylB30cZy4ba1IMRvW0y09kC0KEfVfNsxws9nMoMDjGSTZggXAUhnjtIDzp5hng+Yxw
vDHWR6SiypymDSqwLOMzVG3Cp7IjkKqLGmGD2cqSRLk91MsM9Z387ptPJLX0PeKtnK5SmbGCGAJ2
bidP0bxdYmJwWFW5kgJ8Dlfmbr3puUHcN01fBLBUCBV8F1Rebe9LqAifjga1g0r0xJzW3WPEQPCN
emGCzcHmMFYBoiPKEykt8UYVHGmMvo4u0aVLOCIUQJPDIOXUWXbG8ueRd/5bho//hcp99zZ1CILM
fjqFWr643VhN9OGhjiHFS577YGqF6i4D9f0HqYvtF9bGlynrj0yJdj/SnVDbrtcKEsKhouCJUWSY
NzhcnC6n7QG4BbD4EEZCh+Cnb2KTulWVANrOdS06zCeyVfPUmSkEWK8zVaaHhWgAneSmDU4yytyC
/oHTSfq27C4S7N22FfpetxSE8w1ygHEI7DQ6XpiEvozHMSLcoi2D91jCw5fMxs1Fiod3ASQtaeq+
NivFxEvDh1HxeHk3P6Fj6Kj5LNLBwmKPr1pPWIl6tlVwsA0k9NgH74gUX9fNzB0G0wMdgwIypTi2
srWQTrXOBUmOICh2wcK60tcrP/OzP1u1FVKF5bbY8NgrlCyTZRqUxmkG8uNu9uvQDzuCs+A0deH/
NXeBGq48HCaQkQZ/neeicMr8ubrk2XrxbQ1PGoOFBwOHmcsM9ZwyPZpaPvzccZ3dOm2eY1T2EC/r
Dbirww1+7k9XtKjz7YEYBk/Tq6r3nA7n6W9kHtr3STA/mLrEieyb3GEYPzkXcH/PlJCXwvALq9dZ
1u4um2V4l35i1Enp1Jt1X3PqLDxgpHQfoO3uFUgI73L1QiDh4HRBch++nBrK2oyPSm98RgX6yPpW
oG/6VgHcPetaXWJ5SR4YPt+BYikqYfcHDToMcd5uSSJTLMNMb19Hyus/Gd8pa4nWDuY3bRZGEQ25
GT12GC2JKhzoErrs1PHyAZWPFQ6LIWLEdheQzj2Kr1q+XibTvbhvPczfDyE+Mjj/17eepTDMHRmC
noOrhaVsYwJ5/R5bU/bXgBMZ9UxgfVQN81EH/cMdBDJOSpu9dWtxOSQzmUogYJ7mQV0amtxBoGrp
s0vUYbEcZfmKAzzw9RxYcS5Z2lr0GsSAZAB6U+ZYsH9KZiyFVUXeEujEmWanGsEGnyT/IMk0kjJ7
8Jr3dOJK09aSZVdaB4NCxwvn/UPjaPJ7D82UPh350JfUYyzwEK0bDoMLzoGtwu/AGSolUMz9jtjI
8cqeEVYNOI98bq2kac6UG2sc5NjcC7R1E9bSMrOESCnxSIL8+OczgqgtHxFt2YdJcdUGjNA+RE5s
jQLkrpzFUBwzh2HIT9YOWI0UqV4qDYKMhL5ncGnKx8Y0btRt5oXWuqL0O1DjlpzeKw2THkQo/yAI
dTrdDeQTtaBDowGBklHxkLkAxHz/BgUraYeq5nwneVUlGXVc6JFGxu0iEaSy8s+XVw9YNyrER2lW
BmuQriilfcNoHAY1LyAnXgTpK2/53nP3cxRwIe+Ua/8UmBUTC6H7/hyktLLsdRj8zC5kBH6vtIJX
LAyl4RStZNZubzDR5sMlwBT138YlnBdSVzeu6Y66ahaTtIJlD+723nOCkj562VjJlk1WxEXba8sK
28GMGTh+i7pCvFlQ5920NRq1/vNZ8NYXeGmCqKGdCyFoMggxMELtcaIUgciqrFiPxGcXwrsAFx+2
DrrxXf7R4aYLLF8gPO/hgRpPdBVFvccA6MGG7lAUbRAjkj8v5IOSk24qaAPMwkvWEzc+jbO+Zeul
AQoOewSMbTRlier01NmjAzobRes3Ij5trjmOl9DLBhuEmG9zexe1Qw5KMtjLsPgG0qYtGYA5dEXm
WldfdXRgeBZubvavSjycioIQhOvyOYlV7+6GmjX49xGcuq0OfQ7nYPBlMOnREHwiaOfChRFqcuJ2
iXBFqUMzd0Thn58iSkCX3Ab/zakUjNYunEmHaVn4wXtPxjvr7WsbuUSG+PjlK749jwkgacVwBEEk
+K/VRYB/sJfDtWt83JuLF6FfohlxgzFk3kuOQuN4sLdXi7jDtWjLgFGPkkZqBSKoJLJx6tzzqPQx
0vs+R4eHQlDhTJl/jMiw5t869AvsZqgaDMWtQnW62YmQzL6JUEjdMzQFtMrKSZLh89NiuXDaRHIr
TxMpXkUoaTqs3j5XFqg2yw4WpCsmletY9xnjy+pVdQQc7og7WIdjsmRkVNnOWFLZC3g6m4svoY37
5zmk7YtigV56vp/+YP+AfZ4S7RGUl+0oJ40NqK0UYDnkGm5x51Saf+C4UvcKAa6+Q2nsmZ8KMOK6
846+5+XvQNVyx7gBum6CWFKphhX9X74cRW0M0FlqPi4bjMN87BF1yEVeNpO6VexMPBzrNZ3JgN0D
XAAbSgwhaxyYwHNXJNLto9hSNsOpMctrs/JKvhilGqH3s+bCztlaMruODk87+vkqumEeHXGOYf7t
J3UPXLh0PECEYMeJ+YQRxI8LzgTHsEWwvFek4ORs1B0eQnL1MQBVpDOX7sYaGZxryNumWdVWgHON
zsEVRIfdj5UA9R/fGkk1uL8VRDNKCk5t57+yitArazcydxrMk6BQmhnkeiDr60lhXXsucQ3/23xE
SGzq0gtYP8NGmgmwFlCERvy0AJxcCwAFM0XsSrzJGx3Tx4suzDQVINs7XCiobxXU0f8do9fpg6/f
8KwbkcdUk848QCnzDw+M38fk4/iFcDHpusekuOu8P4bwKZ+z24wNIn/uFiv7Eej5J843JXaAO+jx
1rez45KrCQhYTb9ZJmSfE7vO/lX3KkI76/sBl9DtySXCbrDFwGiBESdr2+BhBDhS/WgtHnK9xPuj
QWpJPrMIqDH3D1r7C+XZ3cjb/078HRDTrEWjBCqyxu+qsfB1+D2eiMJzu65guRY5BEI3FwSelvcG
hTMkP6sF+rGjGVaWCaVGgf/pSgI+V0nIS7cdmyaRGoE6KOFGprqVtKaoIJH7tan00O3wAF0We/11
3Syze9cCopOIAK8g28ut3uiUI2kXFPgbgO19BS43wvuklhmlsJOqrS4pu1Mpr2XKa4MRylE09P2B
jvAUaudMDy4AEIRyGJz5/Ox3nASmcvbkjWxxsE7iEEJuFcfozZ4btK0Ic0po6Ii35HswNHn7IViY
UM8J7iQOijyynwY4lzEZ5m4WTMupIV6HT2BdativABNFsoST69xNQgmPp8qTnOvOjPVGESAL9QXY
nZEBkpf2brTD6VUKLzVg10rL+9s0LulxTb1ivyorLz7rOoCWS+0FRtut2eYya2k4HjnU3TJqZCPK
ee/W49x4G3jSPXdbFBTyrhbBwtm+Cu7BzovowM1JIbd6u6Zr/zgyqqyDXwSxh5dyzQuLS3yiVsWB
SNSjnIL/aJaDkJEsef6yq0NSV2aSpDTN9nnBccKh285HMmCiy3dBNZnXHC1U+q4F0kJ4OGYaqsTw
StaFhuIQcZQ1HuYAs0e9dS3sUQ/jdbz4pcXRX5B/tHv6cKttzwRWgd6K5+K5aikfXUY/AI+4Wnmf
r4EY4runybDpt1jGGRoPkCtk5o17IRKo7Crwe5jKXe4LsxreiB2Owz3PSa4p38htc+OkibNRyMkU
4rWxPNlMFYn6Z/9P9Go3zlZ+qT35u/8rFUArtrJZ4ZfJWtVT1co1AAMEfZoPwhEoHAMpL2961jzg
cFiaXwEWEyw8NUZz3YkGhckEm8XV8uVecfEttE2CSs2aKSL2fyNqoJF+09Hr8D8axQAhRk8XP/9R
RNzKH6R5P24fmZ7dtRgtr0miU+U0lwd9drt98z8gqAtnUe9fKyTQhHBgTIiNW1wGEDoT9WqAXyTS
PtZ+vIISESWECxh2kES6vdh/lQK+i6dc95oA+1sDeIPNPs5jXWeEuaSQoGllGQXxIuZjC9PATqNI
NnZc3gtok87yT19veh/QKcOzVSKuwgW654cxkhgH3/v71XAEw5wlEa4kpmQFhztiwGHETC9Hjkww
mJpORtcOslw4Whj4KOt/8V8/1Mw1TptX/C7zwA3HUJ7ej5VQUNGhN/daZTeU+u1DbbZIGMMDiYcv
WS1uOmhvXwRiLgY2pMCM9o+PaF4ybw01OpY8MvucKu26+LJ/brt3orN4ZreAX+hnDaOyby3I18uS
ReRBqb2U7+OU2tCuBaVBjM7+RPiTIfEVlB5kavVHZO96Q9kLt9Q3EHEKD21x78CGrQzWSv6mGtYY
XVVeYdpZ0BBv9kElT5EUnr+g8YpdCd6M2XSc+RK2WqPyFDSe4CQLwnytMhvol76zKQFGzrgUF/vb
fRmo9hTaEweyFHy/ja+qxJ579EhBg5MixEp5FRfBJhVJDu/Qj1xiTRnA+aQCeJnjtoCxWLSsluKG
6dXMnOMJ2Qh1IWQKYT+dVDs4a91b3paek5bfT4ITEsWaVTD7lIa/19w/9gx0OTJEEKYDO1lUXhax
XlJEhShnyzCzny7Ici6L7NVUbE0LV2U/yOrsbqjZLOaahyRdOHlpCwLgjUCcsm6FhPooJrPEL8PT
HdwFRXdjVdQNdMhBow56INqTbDViEF3H7v7HxlrVgZJsBDx1orCM9k+VSoTe97xxrySp3tO7rAG0
85vE+J6R+YHvMa9zqbZBpT9EVtTyCQ3HhsTiqt1wNJCYmruPJXCxKL/h0YpbhYgNcWVVIMNsMDcS
lwtTEHkPYwLpBF5leOcxf9jJPz2X9pex8DoSY5NivF9Qj/c4v3eCggaWDdxi3cZEDvmMRT9pIdmZ
XJOGEuLNXuBXy4L3IiwDHQZa8Lf7n7+gfvEBusBrXP2IGI2nT3np8RdmKu5taR9QL3g4KayADESq
RdpxAtH+xShXnhUV/TeldduECs5bsC6/4+3kJmVnv5PJ4HIP5jNmNgAalN/4+RnzVqkc0/pXKeyl
3Z2q9/UhHd49mwiTlPefLeiqTI9JSctBXkSmfgiMwaEbiXa1GsgcdRzvgnt4m9uVuEcfcaOSKGYB
EYCam6rPg5XErrwoOcybc7G7OV2qDQWiMwYXxVqxSFQ0ymjxo5JdGlNxmska0I9fvRLpeGPz0IDW
zExqyIgrz5YRuJpyeP9QHcyn8PQ9av9/nI5x/B06u1wXtpjEHBjIMEMG3QeWwa1dTiEtOCssavG+
uoT7ph3hoPW6q4olofFMzGrSVyw+dR1WaGM7H3gQkoUPXtaacvvXTnhx63C5cSMCvIkduzVl/E8c
u8S4I3tFdKcM/ucMUiRHT3sfoGB3N9N5AEZIEUshuM43SpBNEos6CDEZj+KwzIEc4sZWQoihlvd3
zero+wf9AAGCicNGQXFqzrFIfjEtQEcxsK11hh5xraxCP1kBqyXrwdH0OYGgSZNIyqDGCgua4AfV
aVPvbVqzatViLdGjjO/3k+Q+dnVZKl/RkomH7a5p73Da78TrXnM94C8FQjg1IE66tTJs+Y0+Ss6w
dFC2AKV4NAzmK4I4xghuzI0OxYTkEqkJVuATxkehm4wH05EzkKbRpJp7OSgWADtdIaBK4I4Cb31q
b6+hcYbuhds2i+I6t0z852trPUKKEeOyQdo7W7xZz46/Q8//DBE7dg93NT/CBSvUgTZBKuoQ8bfD
3iPp0+ixECYc1uDQaZuHi92g6WbyRu6nd+1r1klP41cbzJfneA7FhmPI/VVBhP8Q631IhQbRNNME
fvPkaKKLiXvnl+FXIUnmSqL8EWjDmgGkKu6rtw3jGSm0nfM5Z991OgdZ74r74uJox95t3Ju8GKZ2
5stuGvu7uYfsOUnbVABOkhJtu657kgQcxowQ5JSoigNXND/HY7B82T5jXjLYJlOaPbzcZQTd36Ob
L6fvHDs88T76tFtVuQBF4tTMIJlLwGnYGG1SQVZJ+DVyKkRM6tBa9u90dyk2x5OOVmTLeyO1jkJd
piAVf1uloRU10oeaDYw2ro1zkn4mZqcUtPSe7NlhSt2PLK0Xv8KD7xEQ/z8yYCjEMK6SFyefepgP
OGMwKn5SRzGWSSAylJOC6lSIGv0E7rvcrm8tvBsNpQmyWhXdzBrRKaIhs4UERgPHdClCnv7CnWto
H51QtjMDYBgbMOmt7r+CjfEygAvH7WTMk51ZNeG8PfMx20T6K/P3An0yIDkagEqnG9vbCTIHj1L2
jDIh68FKKaClYTaA+lH8iaNQUBdWCpR3uPWgPx+gumL5uAA5OZ8escdjQEYXn0MBiQvdB3gjTssB
pgOON9OzXpPmM4lwc+Uzw3phrKTuOc7oTY3OpfX5uluJgGDmdmBycVaXtj/jbyRD8WfwO8sY8Y8g
TbeyCavqWtZs13Aqo/PJzLSIq6gWNIt7NJqD6qKre8+g8T7pgPdJmBLjpH9JmtJidxKpaiIsT/XH
3vFz83M0l2SNJeRnSZh/eCHWFInKLXihcwzVrIxreNJSxPDu4CCBnHr08FB1k5Y82osDB9uWLIXg
VxcNxi8ebz5u5cSYFtDyrIf3NSa2Kom/R9dgrrFOO/BGfUuw7a8XVtzmQaYCXi6b2BUZhozkQUzW
bDaQDcC3FsuPIaycvOOkSa3oKxVplvqorpppp1die3mC0Uu+U20wMiqVr+xktKXl+BtrnkqA6Dy6
7HTVWKvxDJ5YLAmhUcXP2XnU6ss/YvJTziidkp70nWd2b+jCgsiCIJ/iXjIamvEnxmLGn2/cagfE
dINPdURiADDphfttyNmHtgFBZVLGrwyUvXenMqs4vp5DV2oIgq1b26IX8EHV2Vy1SQ74kh2kaO9I
E9jZX0YVTRQJErO2RYeFpt3EtT17rHdzzdIm/EgheGB46QrQqdDQF2FAam+PTFfjO70dU/a4sf/I
/KAk+ZAkMFnPSvw3vc8F8XNMj8ShW8Sqh43SshRwMzktqREBPqZc9jYZfS2wjCUKdrawjXJ/0KKO
yT714KetT3Whp1xXlRjgHpthAnotuGgXWZdkWd7WcpoKRIdFj/raZbtSzwes2+R/vjQWBnbJjhwx
wK8tPeVOCd+noLJVaa8+97nElbCiIlcPuMbt4SwXn7yTW7E26vP6//CloieTjuL/caQezH3C3bAS
LlQDv/acdKhl1EH+1f0b7tKviVFkdk5qFqBM82ZuNSYUQQJnJ1WxrFprSQK4N3yD1Qan2Jf0tsK5
FPHtNPLFDQwKYCWrvk7IO81dy1Ca1/9+6xyo7I0DKVlW81vRkItr425DafKw3TgrN6Vv3N0I8xV9
1Qt/rFW7As0E2v+vJ+PkNixFj7sR3XwLkN+kabVRLrX0uKiCsaa+2/H+MZx3GnP8cVHWzeM/n3Qq
YBbVPWR04r6fohXYfuh4tXWhm8Y/0k/UI7if6A1plmI3rr+iYr9KiJ8i1ydNnv5zkEiwcVH7L1Dk
8mlQr+Pto6OLkXSJwDf0foFQDedsVxWSFCskvp9csXwzuWkma1QsflQYakmBWZUbG3UJwWnjfNGI
g3KwEE9ufbX4PVUbYdHLs3dF4uK5W0XzE+CGfnxOlxIJs5ZQl7WbH7jIDPJbz1g4XqM2vFQFtRvH
HyKbb1U7H7PRPQwvtdbpf042LhLdDOlk8gruIlob1m2reisdzF4GG9vyj3cFyi01aFQwJVS4z8QE
QEa+0Az/HkMm9CXMQ1p8zXBOpwqiUkFTBmB0INMyhnWswLPtHlDqEPN3flpCZxAzmY9OHH6oQf71
CUtcfqN4j95tuJ6Mlto0cQwUHVNHyrFOIldPFYA2Ij9uKb7cA1MVSdLalIBkxV+nlqK7lAQb5kLj
IvdtuYHGXD096mHL2NzXG6mNBWgAY4AQsd+0KRzOLeOcVVkaXW+wqMlhqoAuNTKQ3vnJyEAMOBcx
XB78EWGohLDGgkEkXlnTyZehQttLl2GKsFWzDxhy76YkzUm3G2EXcoZ0v8rQ6Cu54ab2Gff0nFvX
MKFQmvsMHGuLt5R6wO2mLfaX69W68Aj9/I6sUJrQqknbx47oFlVv671lyBC4nbIlkUsUcxRCeXh2
3O2KjelK3JOxFusH7MnxDm8F41yU7JUFjCdAxLpKFKzlKGmPd0XnEOO4iTsaVuahH03i5ITRINpo
atEIBetGPSscoLEsjGVQAC68tefQXUwkjdgLTbc/iTR+PRySOM9+S0JPNZdT+YqephhquKfOSjgP
sViXQAuPc0vqWMbF2BWqpGon353ZYMrBhY7p0zKbvPU5ihBpZKRDB+3mEadCvr/V47tTxY8cPwM0
EZ9NzMWhb9UmB6aXQLoG65F+BqsY0zujrnX2M7hSRZ2bLKnW/cxTwcz9vrhVi3j3zxlAv1TJyjyX
Dv+iXvk0wP/95lgqBQBdxfbD10v+Iiazifb1A+8KASjs02rYB1dq9FKTS2bOK0GDDSJ49Mml5KL3
vYIb4XakMEJIHQNVbE8M87FZpBcdVGyK9OxVOFLXQUs7UruH83hq29SHXBcWJLisWSWLySWpDFB7
qZqNT3EDgG83wpRLFd3BZlU+/qO4yliByf1gE9MyAwx9OKOgqFsRA6KHMvOJ2/bVeveMKl31shl4
T1URFjmP9LvkeqAWm+ZKwj+aSIi6Ul3suM5yf97VssyMIAfW1YhBe4FZZomsTOLzmXVa833+dGPo
kjpeX1cYEStpcJYgZwWsMKPPYXQ0cebj3CqJciywFt58tl3D7J4nenXHQAI4/4shsA5uUlgLSFbj
XprILzYlkyz2hH/lMi60dOQodkfNmyw4/AsnIRrTsu+VsMa8mbXPtMxCntF+7i3tEhq3fnfBjsIB
PahKMF7x4iEXu1VDHHHRNfrj7wLZy8KmPBfUm6j9VB2Yk8uQqlvU83ZkP23j2adgDvjncpTfufiO
Rc78SZyaHNDlqZstUGhql5z8WRH07yOQsQKJVUeh/lpMfviHXRSRNEzDrTU7z+MbY5L7N/rI9Mkn
Vb/a5Eh7zj7F4SHX0AyFCQAAXfXHW+90b/v661sSvjrhpquf+FWc5ozGthq2W7mXEF6wnmd8ZCwV
Kv65oEllJ5kkalAlrZpvYlzTWv0OrjPqzuJ0Xrb6Jtg8fFFyKljkYmVBObaVqVqOWk2jQ/5WFFZY
Pm+DOMH+NCXtCTRHe/CCNp56hlAP32IYty3MXAAGn5RO3d3EZQwnXp5oyF7dHVcSEgvcoSspPEJ2
tz2992wGJ9Sce+Yeou3neMBfvKaOdK8G4Nb1deqhMP+4lOODBqKfWaOXta/2RRKrggNWhQPkXQWs
CEp/oUglEEsUAPtXJgDSXFLrcLJw7IPubE/00VyrNWd07sc5nktaLPANRbSlTdrlsUOOQwIPq8Hm
fL8mPoHxbRdqDKomq/S85/TC2o7+5kQOl5LxE+WsH9WzDQWV4Ocw3voVmatpsKY1yekrfsf+8xDO
2RjWpO9CIvix7SsE8YSNneKGXT+9Qz5Rty0/bEIJd9XgnDjvC6WC4hOvDCpBzhHI9g9E03KjHhje
f7wUa8fzUF0OgEwR7iw+Zy7vADfqR4gLxqQaMSYkhRqzef3zEbxe6k5NX9gyb/c559zxiTGrd8gy
AQZInboWx7I28Bee4oRo5s99mXUVl5q7Wn1QWVw5k2E/k+ksZJMlk2VncDvWS0D4OlXKnyN6ZFfy
+JesPv8kWhwZNynOjItR259lkkFushj3WiJ332ylC3K59TXYUacXBcIr+I8Mwe7Z25cOy9MZiIXs
jSOQONYErzABbkJB54SNhWhqS3msIsggNx7iTptei4WIEafLJG+Yyf7SdkHiLXtI9c4gdh5Iwc7V
Vc8eTTB68YQZRJLvyRiDC2G4JJUnT6qVXSyfe9tX0tyoT/VizDaUEgY+HSmq05RH9KZgvwWghmYL
i5lodfRngNs44Ydh3h5gCcxQGUw/jadMah6Zq6CMYVeqq511JOr+e+7SeCHuzJKXW4g/Nn51I3em
UuXwbKPB5p697eLtWp4Ii0inqiuQVRo+z5yRItMCR4E03R/BuJRbi8OqrSxRkk9SQ0fSuiN8lT6a
YI57AGcB8hqZ1lnRJGwTZ1DOrQXUo9pV3n+YUprIMn3/ZnBa3F4t44BYlaSL9+8XhVcyG+XDVp4t
qtZXm70bXWB0AutEFL/1YO6z6Xk5547gaQt3EwstJ6SlYJuRFzkHddU6NfbfXhPjLDN0SE8yBbZD
E7yMgiLgBJTY4FuIXIfl7JIphsONh2k54Q37oh+n3xhZ33lYd0lHPBEjJEvdF0MXPpFtF3/8koVn
mQlXmjRdo3zVkr0uKgTM999fEK6O0ERp0e3qGfb6hJmz5gmMPIVNcnGsoUcCrfGGtkWpPgAa0wcu
vlMMnv55CN3hLbEYz4l3gWSugWJHTjcwRwl8Ch3YAZvMIwFoRegLc0UOrcviM2KQqNhZqL0CKpMl
sSHChh1FPl0kuZVSFCCv+YpbqloaJEr+zIIB43QWOCCpNmcUU4CY4Wn7jteIAlDygRsiF5LyRy+s
+SOeIfur1cgotCsJdCig3fJTf2n4Dg/yPjbOiD469VtuBeH29n6dtbHqZpy7jL1VsGSQRSXCmY2R
z+7GIelBmtCM6kOCIgJJpi01/Hj5CqLryx4Kul2E2omj3XKn9g+f0lRgot+La3F0/HGwfgcqq+47
CcbLYXi9A00wC2SjbAyI21x5MW2mwfyixgiBeMNWsp/LTl1vZ1eVEkkI11D21kT6d+peo5ra1y2x
3VxSlYsl1MdaIJyBswSLfzQv5l+fgPydoIaVJJvbEaSNjL8d/+3qyC8+W6hPgEhWZTPIXCNpCOhg
ZlX8OfnusD6JWhOLjyHZgOogq2n4jxDo78ZqnxGTeT/nY/yUbVgSKPEqYbLnfMZTvgQ3/ID7ox8d
ru2Nn21mvjnazvnJnEKiw1LTQjZQhvy9OiPlev+o9H8afLVZp8hKCpaNoNnQlya36JCqaBuEe2vS
4azi0bv3cAfWwDStMuqvtRbgKduiRP2+lXn57ghAgpUs0pN5ofifWQhMYc7k2ntRkZzB5J94vmsz
bMOVvempgzKvflFnrBUMB3q7ckIqU/0zzmFMGG+wNVKIzNeiN0siGJsUwvWu07+6DEMLdZADR37B
G61FbwqFOa5iDCwPQKsl3jSXSvc0jEBKDrJlGl59XclS7Kvv6cZfKRwiGOhol99X6ZRb3rD2pN0L
62zU4Z/+HsCIPgbzQFG8FCNUbMpIBkIQvZzf+4c2kcKS8AIa+Y8eu11KctJ6TvQTnLJ65xQCrg97
kqqKfQleaWOmrhzki3cD21Odm/ShWiZ/Nw5Ja99i1KYYxIK5lBQKpe6P+Lid1VIaHrzL15e3Th49
BxONKJsSWQBQ24SW+3z12JTYcBDW++9LZM1UdxeWRfVoLNftTxcu0aTV+3ltKe8VFcD4kbpGmBNy
7lweWz7Q/bxUtHjAAkbc8E2pRLe5cjuSTNki1dCCemeyiBm0wSBlCxB5kWySe88YUBFvK4zkP6f1
jjyxGgCPv4D8hgAigdP6hej4vToJLiEaWmJzBwWfdidgDQp91WURLOyWE0wiEG3T1TvJ6GYJl1RI
vBxkNrHlQkadQB1yUOezn+6J7e8NEA5V1HHZsJ+jBEqLkpLf56+xHMBFMFG2+aUKMBLHRrJNCCIJ
skTH42CIt8WcQhYxzTp9SnH4pWjm0Qb88DvJ7f8WeKACiaiyunjmUjw5ySsr2F08hKslokRjkUo7
nGjoeCdMwbCM/Z+UBHF8EoB47CoVZPChwjHO8ta3EjLOlHtUgDgyGLpit9ZlxVLr+j1dJcWvgIHj
ZZBzcdqxKJZbRnHvdLt7+5uWrrH22WU0Lglb9coiXWNXbT9LAyX11vIF+9+JFGKssYucXzfCa3P7
y+rLVqE5NC0vK9hYhRNr6jeeVFc+IpjYWAchZtGP/V17SZ4/cu0iIyRbRTFbEnqhkYZFKn7Vhmcb
UTfKXJm5C6st5C6sK4ObAi9QAyVzUGTk8r26ESvkhcn0x01S9jRSOfWyLVrZqLy0iRPEp52cp+Sb
3YfgTn8uXmNWMsFTDUWgQg3feKkuzO8FdfBkscjSLxM4vmUUkApdaxK5qzBZa+hdmlV1eJaV0c2+
WD7uzWY98+gtiORu+PAZwXGSSAgGg7R2nTy3LzhTqXOynqIxVedvPPcmr/yxw3XblwYy1+KhSEX/
lRipfwdw01LqF+Bzq2/wnqwzy+45TTN7hQDExlJE3RJhDIWO9I+T1epXdDEmToC8BvoXu3RsX2D0
x78L1dRiOyXobq0ikkBHrHQ2HZkJFqN1QXS/GRi2WN8N9einZEMfcQB2aFy8ZjMDbVIMklS/AYsd
+XX6sL9AgThxMrHVcZWnOGX4V8dlRt2HbrEcL3ogl25n3OYLP8cUJxxAcPDg6qiWVpoojZBJyoIR
DhzPIm/vE4FTG1IYtHAAApg9GUTc7K3KtyDNDtZ82WWLSwQEgYnvk2WUcoigIju7HQrftgygJlFB
cVRa4E+/4gzlYMUDqZaSLAU+H/6aOTXaGccGoPlIunVxlGC69sY2C69WKT5Nw/RAqdWp3ht9NagR
qL0dU5sj2+sfNkn5AgE8yxHp5HXr3dckrH50IJs9RAh39k8V+zpV8bEhbCRankBtfwXUc/IG2h7A
RSMOMdig8tvZPm4TfLZ0zx9tvQy3jBSVPcV3Od2ZY1EoGM8ef04nqX2MAl+B7r/59wwp5+M5Ih0R
hjlGgpyhKZ15zijemp0btVYyVstwuhVjXVpX5tZ1xO12f6fmxnXoisQx3wzaW1CeRzMAymtE8SDX
6jP60P9m1882SBYXIHSkw3VJv/+R+ZKLGIRk2iVJYu88HSukB6Qi4R1Z/QYNWAiL421QjJE1sxv4
74W4h9G1y9bm3et+dC9feuq/cW7J7DW58r1FeEzBZ1cmupveoQuGsbJKDJm8OfVEgIwDjFl3AhJa
yG/i+0taXtIGn1q51/FFYylLmIl8i/sk12EUqoYBXddcyRfbrAB5I5GcYgfVV03QXTEE5KyB1ooi
KbvCpBKqIvw1mpbHuiUfwLwRbfCRXdUOli8pSHNEYwmAm4gA6ExefGIn9oE4iwp/nJ0MdVCNxuUt
/VpSK1QD1UlvJ/TrFSboaabOpcRvU81GF/3Ljuym+RdEP0f6NLnpQCaKDwGWqQYTn1yMdwMK0OcP
eOEl+7pe4d3KAMl/eSVtAttfXGLKcM8QS7/G6mQbNaVdLT4wibB3BsORAWK5tzEQry8tymiUGtwK
x81kGcFVShBTQmvCgZDoFhFRhcdaikaYqZUK4ya4TwapFZsrVYne2w/ftn4Zg0vrEob85I99eFNM
+RxwZ9+bdAKhWbfr8+xvn4Zz2S8V1cu3Yn4cYNs8OrxVbMGCHuGT6ZJGcIiP65+tTchYWyybB0Av
gR6wxCFcy9NdrgxGB8DOYNDoWWgWylH0JnGDt0r0u2WKlpO8v7Haxv/wXhIZ+VaxsI/mbdv+bJxI
7AUIzlm9CV7/X8+ECjWrvcT4nSd9cSC5T9h5rAK8hnbdY9XH3wlDfZsAoA+ePLJkzu30UhLWRl9e
vrSr4mopQUwzZgscv3LfpVA6b/0dRQNTbn6g2+SOJThUX0FUbEy6WzuG2UAJJTVDn77pestoHwsR
HuQI1Bs9hYrMEh0bMELtmswVb9VxldQgJBfzz1oUUUfRkrdvdm20Ss+kmaczHfjO1XzoRdt7xnrg
VnutJj0Qw4EfC8KfhBRWYbe6yXyI8sHQ1E3eSIAF996sIYZmzWVkcmH3A6Byz5JBgO1KW9Chc/xB
s5GC35mLWVktyA2Xk5GNHYoQW3RWEseod99rHQyUmdNnTNQl7Jve97rvSltAOFkjbSvnLSeeCFUY
MufDbiqjWubWFnaxP4eLw3Qwo2VLbjN0DN0t8I6PhpvOQ1LKy8BO8qUa+y4L0fgcecOpBlqriVOJ
uG39x4pBzFzu9yXmCec2BOtysfVKyeCy19/m3oTAqQshxvWM086z60vXo+MoCmsS0YY9/GQs8Xno
n6HjsUp1eqXBw5kkN9gbaDP7aOih+4nSBeiwDMITibzGVQx9F1+gVdKT1KE8QTuqK9DF/27BNEff
gemgAFW6aBMZRsmH0uwUU1R5a9g6G2l/Z2tmyNyiIOqA/0Su2NC9FMmYxyR/carAyF3M0lj5fuN4
G5hED8eayucE4M/UTImOm/Og318tQ0Z6J/EiU9y8T+wSnikKug/Nf4GDr4XQl2ZdYI3vvXxkfOnv
tAFQuNVTiPsPe2ibzshAzw8vfUpZrYVywEJOMfyffwbknuE7/w/PvGfWEZgWtfkqIYJxbN91SYqM
Ss4pJhh7LRdkcLFMitERdiVzRXOoEFCvE5ZIwolL92yov5B44XvSgRkuc3HT5d+6/pK3ipYb7Dzs
IsWxJIcejJwsHK4SskSOyhmK1UECvprVGWdYFl3BNXhZ9yBgx+HyLweYLyGpm5sDf/8EeqfzL4Ci
mhCFqYK50gRdEuZx5Vym7t4sOdc1XG77N32+fmixWt64ponHDtFgOkv+Pn9Bsk088hvVYhc5PMrB
t1+pMVKFk/XLz79JWjz2pRYFwF+r5xhXqDOkF/YorZZ5KScL5MIJNSnLC+VzimgOVR8EOqk7IyfR
25I8cdHWjp8VKRh5/R+Q3q+EPo3A1sEuSx6rs/L70lGNATgymTsKVDwZLgOudzVgpe+TRq+tdvww
4qlqMsXATnhcMM14hJXoU2LOLQpAL5nOSetcrFNwUaN0R4GaukwR3cKfGTFKMH+UYc34g+vSZddQ
PT+n23pS+lEjKyXSolFyNaNQfGhoGbHRNJH3jPP42LZ3kj1LAxDJoTSr7xmrfeBXQzjtpYZXNOkB
xvseW+jWQCD0mABSpfJgkpZw+HyH+LV+4enPM0OCowk79Zs0CR7LZfvRQliWwd+STVWsL8Wq3j6I
8VlAslTaXlnTCnGApgqhnLRGKmMIhGL6O8LeFo+frKqsygDTR+Isy99XRL+KoMRhhVnJJ9+eDGyd
lbh8ZO7wChmAfXSk36ZInglsXtcM2LpzKcLtwVNe43ake28GyLdvZDv+P9ihKdr9QYaRahoQS7pE
SBEkRSe/nbzDTfxx6kpfERSZPwamVvN1t0e2xS9sY0xq2oMBnYIK0RlQR462tU4Kwi8ZuieYheub
19dI6i2/ap/FF3mqtqCgLpeseVVQ8KFgz2vVyBSdzpS7WfdfbZFpKaoJZMFCGVLtU8H5J9oMdQmF
I8MrBPh7NK+vCYYbUeMrKrJ+oeJ8ADY3MluQmcvj1s1nuzAtraw4Lek1sW2QJqU3212xvztDI9DL
zsp8lmn4gYprHlccM+jSs5ZnPKINKp+pZE/d7Fv5AX9QlufzpnnM2wjsAof/a9yeQ9KO34X6AFen
r/pQZD/IRBfuoAD/gkl3EwK0xV14gC4dw+0M9sSAcBxNz25gUVHIHv/U8/KKZfRO3NgAPUfNJZys
iKgWV5n20RWoRoiSxzi6VDukqyDikIstngk/8ZFahnzImd7CgCr3B3dSwd66Y3RKTM+0DlxxZjEk
AUHdhpyuQE2aGbg4uUepUuqQm8YPTG8xj6VExdzokR9xCZXxOgrgKdB5gvyQa6OvIiRmQUMam9ix
pbzAEsxUjuXK/lVPg877x4rJacSbPXf6Scpt3z0xgrSVb+TRWxMTE1gk9TtFFx8P04B3jkcxEwKP
UyxABWf8SdjWfg9OUzS7G0JEYdMUqTo+zFFqzWGda7DY5ynzoXzHTccuY13okIPjdgz/f8xl6GAo
PppkabLo983O3dUe+uW+7qLzdahx/2/5BQPZ6ENOMts5qFWGpWQAZLt4aPddadcyZTrLVd6EafNQ
o0vhj4S+oI6AUKNIXgHF8cCgSVLosIABKYGcJKQV+nu6SskBwpVsOTEM4kVUpa0QXmfDcBiEoB1o
bHbFb4V/0+Fg8oEo/o4/daaZVqiiONznRvJPhA+Dz6y57vZPG0MqHklFTlNomYcJM/tBfLdT6Tao
qM9sCVlhYEb6RIEXceHVI1ZN/iqR3nC99dAnKRkBoW7JMyjDkUBKXlNyB1Mj5syHduOi/+23octS
DGX1Tnb+adhud28QpfmXu5AVkdkweGzcMkKq30mbIMNSEuTU47GwMX94w9KopJs4FIlLgnX1hVjk
YxwRDgkraNPb/rSaAgtSD8vUfatBcR4jV6kputPypRkjYi/UPK0xi129TBgWj07n3c6O0XmiCkL1
cQ5L2fdC6p1+4qmf9m28Doy8Gtxu3hLvNH9wevLWsMbfeCC34ArH+dZyoz/QBgdR8VOBkI4EfJ/0
2Os0+8Xqh611Ac45CjaC66vKqhoISortjk3XeD0CRwjh26T+k3sfwT4we3Y7LUaD7Xgb2wuUYHtT
YOEB+qBuN7vgXz22h0fkp/UkFh/zLqJZklnJ2bsAYENmlWkl4ovKeOix2FQLysIVtPXuFlUcLaoo
ewcGo5zeHszyGgvYFbWGrbAX/luPymS6ABw244MTkTEEvH3XddLLzL4itN9DUeSLJKFO9XhjSwru
yexJI3SRHpP4KSIUb77gE+YV62TJ6qabEU3HROch600r03pLXLL31yGhX/JUfcP75NbLL2xNhxv+
RZl0VwR+9zUveFkyzT0YC+vkgWctphdGQgwqfKQvv9S4EeKebTCspUc2wSXtzOMT1amZpk6yHss3
x7nznwv5X31WmME3s5D5ZqVcn4xR/8J4yFMCeLmsp8Ieq7KpWG6FzdakCoRcsniHNn8DyDLYcowp
RVmXW69RWZRVTymUZsBkZZ15K3dNCEjztJdmqSGzBDAYuz8Q7HKmMvYGXRXgER8JfU9VvoruRqxW
gQyDVEWWbmUgSyDd4xroiEfCsioIPsbiWs+WW7V2a8i1KsMWcdGCAg2mon8teP6xWi11q6aI0WDu
uJyoJFuikyUpBmONzhSllEvoKTDbdbRuvuEI5gAXFLbF9PX1ve347xFAfDn2ELxGYfJ4C+umQ6H3
qJ1rvKQme7Jc2uy7/qLT7/b/r7757WJ8tGcLea/vgyfHbcBjsgRqfo30XoOlsvCiK0XPhiSBRWRN
06Zned3hqzBFTIuM9bcMvLrsMHhGmjGXgTazs/XVeRUgxl/L1O5m8oG8qb/PwfdeQHve02c3FbjS
qSvA5RmRXRaGuoid4J8LkzJ47eWQSjaB2JDT/P/3jvlYu+P14IjITTzdp7K28BNupmQYCNIMQFXW
MbMPxu+avt2rqKVIXYR271D8zxELTJeHaBcrY2vmigQUaboG3GJYlZISxASGrKEC0FPZUyg9Z2WV
D3d4yALBsSWmocbvsqHbfWUZXY988I+QtTQGV45hIoDpp2uVxSClxDFI4eDpB9hYlz/2KOBCqHPq
xkhrCQT/Fe6BmDPCJjtbFZby5gLIXvHVl91KAq7Sa0gkf5KLFMHXVkgQ8391/nBFZhw55QP9WZKa
9vUE8tHnH+JdPwSTuxIAdVtDpvIyhyVRohfPZZQzK8CeLn9s2o9HKWLqyNUiWGvfgUJ+Xn21USUZ
DowIwvoyr1UY4lGq0ZWN5dcqNrsYQ+SMbAnwdj+Yh/wHzpY1Nj/ngC/J9PqvHHVleMnoQq+5wXr9
RJgdFqDhlPwfLoRuVsAacl/MrOecO3GbfiHLK031BjsgYHcMaQeVBPh1ZGTShJOnbWvm7IS8MTRD
wytEvYhqk+tJCjVxLu5WrAC4dt5bcFHjAvpUBdxzzDhbTh8vh4zCE6jHH7nNRw7vXYakgF9ZwFxO
H7xscDBXreIrtstNVR3sB2Dzc1YnB3BVZXfoLrT8+NeEEQqIU1yydQawh6n0cpExbOx3KgW56EHR
QrEY69ZXPRgU58RiOgdw9WqrtcEF+Ncdp4SwK+O/JqK9gfmBdWsKcn0L5C7uLxZSe9rhcday6cwl
GZIay4uvbDOiP7VD0Ba88PFt82wLizm4h2iTQJwW2swv9wlH+3cdgaCXhl9IhXhV9ruj9ZbM+r55
WS0mabDbhu7r/5lAJwJ4niR9E/CTIUylhBGPdMMVDgLWlqjjFS0ya4PLwLzOOAQ2hi36Ffd89FzW
Qhpiql6f0sQKnUIUuJ9S1RrU3FVLT57avkDVU4xSRKfe+uStcqiDYuccsFvSIlGZ475XVESeF5O0
aGcWabymlLE9Fz0Ue2sm79qOrudiM0NYVYcaOppf3RxrzjJKPKIvqV5xWIHXZJ5PX5PYJXBDi57K
5K3/on1bia+j7QtMU760+VJ6b6AQMXn0Uz0kSEuB/In0nFes8oBIrFo8WNj5NsEv1Kw/QiB95rIL
/GAl1qzpkM0Lw0TYRxXxRDl87QjxIxKVtbgY29sp4kdEUcAlDHIpSw4z5HuyS69pSSv2v8AmkcES
nc4/GEPRY7hJFcYw/kS5yWttvJvdYPI9n/fBMT1CvKW1ABa5pw+pDcB+tZn5YWw74tOhPCaO/ls3
nFPytFeD8cbc2fwAXriMEm+Ne5ONZdwFM/fGpEcNtKsm89qttyRRFzAIgvSa7CrybsAXzIBkqUK2
cRb6LFHJ3gE8KJzEpnvb80oNekuiHVqdi7uHW/Fb+0/ojzNistfAY08Y/qA+rTHy4rEaDV3Jut8x
ahMEGEyoFaC+l74PLogew2f+W6Vx/PZxwyCwepNXxH+OInbalsWyU2YrllghSfe9HTY2w4LI1g4a
HgP0oA7IZMugygN5lc3/LjmlPYz+u+bjPGqzrMd1xFdGGLd2iDPOF+qJSThjLlrpQIg8H4T89Lpg
ZBHldJMMZC2fVnUhGhYuZks97wQM3V+tdaWF89Wfuapf0jWoHRSumWn5KFHEAzMQxyfDub/2VCLv
JPNaN4tLCrEd3sfcdUOan4frI14SPs48xultTLhYeVUaOoHTuBdP1ZbIWaJDzFrRrdlYu63LJnS6
CbYKZtu+e9bo9LIcOxNgNhYX+vjHnDIiJ1YdmXvcFs/scyzR4/9ZBxhT8A3BLTTh4Z1l29gnxlN1
hhUlw0qVPyRkyai2FLrIi1mbxsDalENkNGzowSnNtVN4mHP8CCzL8XGN6wxZgm/yfg7lxKf9Bz7F
C7C2nYALILOTYwRGbxA6vpcz5gcMxCVRuymdLvzaBKVDgv/q8dApE5nLL25AMuawRNZlZBGOqinx
pTs8otbifqECAIjBx8S8Lta3g8NtSgAOpNCdgckrU1wtW9jWFumVifmUW9DDGYIc7RKvPnmJgM5L
CYRujFd18Zy+7XK7LuIDBgigZiZXdtG3a5aHtCk55hVCkzE7C+TyYcqeBsIZk32ETL7WWlAGbdrM
YoUc3UjfwtcoVs1N0gf8dZAVHL1nfjFKHgmYXtiTtqUY+n96hcm74FJaaQNCNbgBFTgviQS2rzHn
+vW3ZIPafwTcTCbTJ9C+zKcsQReWQ+2aFh2a2VJOYXf06GGmrV1Htf0rCFV/krQvuF6CKnlpaBUZ
cpeNzl6LEcO7h7aMF1yDqRK3xBPFAU7bT8POzsWa3Fh2OE9PY/NtSFSTuGy8OiD3eooqQFFHtXpr
QcW5/9gfkkVGN2I4Jc7ypj8CklPhuyGW+40flLqp/I7BS2+LFgG1xvIfRehn5cJJpEbPoYoz3ZvI
H7DMHrvcSB+9+twQ7eb2AvgqU4wflF2PxKFiTvl/L+urHpJ+3E/8QGM0mLEfqFp1wrzFWrIeN9tv
QVCuhpg8KMk+yYYh3IozFPVPEmU/jsjYBjByXZ3eJ2SVq3moLCp3Ij72nmVt4OXWKwBISybtqdSP
8ayeyF5+eJIxl98mJzZSvddmX5f01Vo89K1+g13p8gYRtzrNmaNh51PlZpFmH/aV4seBHT2PNJnP
zudaRZug1DpbK34L9Q1bvW2nav5KnzWSv4dhkVAop83npor4K81akvQi368Y1tF15cYVtr/5Mlso
p4Nvtg1EoXa574qHmWCyZXcgrmjcczIEvxbsEBtHKQFttH0YGf2NPMzt0gd15F2QvlxF0nYdGb9t
YT1S48Zj9KzWsCr7xNKdw52GxkQZtIo9XD2OU+mzGoh3MVO7rSDPNgakGzTnWQT7vKp5szN9lXDX
9BZpnKJ+WFsjPH1u+kv+8Xmq9XpNl5ZClTShHR7xQLiJivi9lZYc2uz3b7ouD6AQ3VHL0Z0gjzzT
b1A3zUFHl4wXTwhbPwmUw7VAx6oHtqxCKkT5nzHlXJkeK2cOiUtEGfUYQgZsbzJqTsChjx2QBiwO
xIw1PiM4DKvSlYwIFlgy2zlz1G9qYLGszfmBb4fbJQdWQNpv89Zpye4OWGQqriv76COS2UpyUO7n
bbMWakIRNlLQAJOni4o40SFINgv6J3102MIggSgYoBPqmW+Sui6OIaJfj/ojGwGw3tIe1aElRjAp
5GuvZMYT9lK5E7kp8m1e1WDzMu8gaz1tXmqpiD4pM9zrgWaxmO1WBdlDc3zj47LCVIZNCreYqi/a
BRVgC3E+tlJHmaX/px0Rkmy3+AOI+uiCqf8xr8dwgoBaoEU8MB3GCUbzkwUuYHClcM8/gj1PVwYB
FJOZkT+dQJ9pmZzOKq9z9ihRslulO3GDRf+ZnDPbjxKGC+nSFyukwoWWXo4ERWpMiY8D1zGW0Giy
IxBh1OpQUBhJnqXHm8JzfGoVyq3+uc3Qj+FSGPPmEVMhdzO2Xi2q9QcK+ZGZLTX2WAFvTQnh0XTI
97o1IOUJSRZwck+yjioJac0q6MvywnnETCi0W9hPAzPYvT0S8E+7ISAmuy7OJbUogh2/kCJAMJ+j
XbWfz2RVxzGMV42njCo5rXU3ZAX/XDPB78S4XAPEgKn8Kc6FGD4IHOavA+YO4PzC/6kb+kjdvHev
PQKEFHAZiPBbsQOmM2phPGeC1kf2LDRq+JuKgC0FxgY3W2ChCcYWi9nwFUfDbzIbxzF1S0s7a33b
IwiBjhY4e/3LJGH3iCz2IscR6+IYizrcPKsK2NU3Je90oEc57fJHi/r3dwpxw+Z8qErfMvZ6/ye6
A9evW4z9VG6laL50Cox16abvZRIrVwX4qsYMcnZEXsnzDjBh6MhADvcJG/bStF3blN6Bj0djXTDS
x7aXB/OCVt+MZ22gn/qfHRnUO71YHFKypsDLxtb9cz5euwSwb8bLGqTdaWJn+GioXQxuwof8bF6/
IX2K7wZQ41Y3ZvGB0ob/LgYeO8lNkumFgXU/1fO9I4o8TY7F94LwNz34g17LtG7HsJuxJwt2SkDW
QLKlv+0wrZcXHbtJFCAtgRvV4DG0sE0VUkXgvCvQSbCdeAho6QyBepS/dbs9jFfqcBipfgp8vdcV
4bW4z0Y+dBuOAqH4K2a3Ah3xD4gaKY1vClcOW3K2+KgJr0jWU45FtHxNutHVz3Cv+eqBHYEUExEC
9yBM8J4AEs80RM4/kWg5RKuManFRiDPSSsDQ6uenG+pcnu8Lke1SLK5IkQTgyEjGiF6a28IOgF3w
W+l+FZJo8e3cItjVWmC7GzAeisMG2G3YqaYkDXbDzoa8x+Mun1/tdw+zItU23P+RUhf81x4+XV9A
NA/AevlAeIFSCw04BDf7P0HC+OCuszVz8LFR+EwCvzyGOc/zxeAm9a+eXQGt6keYTFdIlOBT5T8v
0oFv0VQ2PuTtq/EVYCi2NmKLGvEJ4mZ0KV0CwdC/JyCU/7f/nC0XU404dTkaXbMFIGVEFOtdFSqr
fl2YIfZP3Yh6BWWbhuoZVsaVqljZdE/T1KonmuGle/RRoqkhC0sTJLrBrdyaxSQhP/bNx+/vXJlu
h1qWZh/HeNXWBD+7J0qW5e1O3lmt1fNtelVoHuCQmGh1XvozTpWcIIhyX6dOFzfTkbt9lpLgPNt/
aSDV1rPWz59zpKw3C5rMj3khyYD07n5ZT+foRZy3P6KrF6UyrbcpuYv27dlPEyjPFcg2F9dXlzWq
H+8KoDA7oQ3x5NFBINAb4ri4ChmDi5F3n3eaFzoBDRaFoTz9E0mju9hgSru1ycEYpKUKPtzx/hHJ
5cBloQbth3Gf/euU30WlWYeeKe5SL1Zxf+Vr3wps9JpOt95au7ZQw8ytFhyuhFJjydfd3evrO3HR
9cH681BNC+4tCQzjqvl3IvwelO32PMJwPw9CvR1z9gl1WHJf/XkBxvPLib1sk7AofzEq1VaJWYkQ
FQGqRj4kZWnVns6xgEVgBGKcJArtQww4Je7hiJ2t+QjadJOKCRYw6Pm52GClJa75XxOjHfMS+is9
9F8M/7S9P2qj4d+2q2cJU0Na5FlCNCZC4X+RZ1xmvYIr9Ar0MeDCZzjvCN2IIA0XIO35SNmGu/xB
BCOjsq5NtGxh8F0r36g4NRGsvPdjdH06/F3ovW0Jg/pGKYji227h6L+jvuLUJBdyoB1ICNJ6YcL+
OoJv+KaUnka1Dw3sScBtN9y/8Q8cJXQanMt/hCxc45K5BKy+3dGXaYJHGJkLTFrHPg3en3NdiT0E
QyKZG90xuzmRBElfDT5HZ64oG3968zsnFRrnVMzTFN2hkmdC9fUBcuU2VAm3ooAa49Oq8WUUBJWP
Ps79Ix+f7R3CfUufsAC9IZTUDWfQELyCgF6WYcBGVcy7GUh3xLESt+xGgGx3cYlABZ+hi5VIcgTd
4W7chU/YUE1ONsWbr5AMv0Htc+788aZ5Wab51+ZUKOGJmGGUhW+6jPjFu24DVc45BJHHeUOFAOZz
//LeFPcq9OO+2voNAFZfEFpNCJ0spYcyuRt8ExcGWEtHuoBa5TmjtIRlz+Q+jPJKeGChAkoHHNqn
1Q1f+PZsFvjV+ns+o0/howpE9ZJAVyn7IidmxxbmibeszxW5RH2f66a8AssNn+TE0cG0abDxB0nr
/if19r9vbZBhA5g3LClliBnbDJQLbzL8FpWer9JmZY6grMGpl6j6EQXcp1ClR4Cd7n++7E9lJNqz
HAYTmGTw4DP0ycUDp78oz8AGB8X/jCxoVAQnr4/oECrbLIihNsSC9r2gb8rST5AUhI23ToloN//q
MsbrtdY7469Xf2WAmxzlQ/WHJ9YGxyX0KOycQxoxSqgxssGf8ClnsQcTKp+L6GP4pYx30yb3CDh6
hMHBAzKrhndqG8e1gfvur96wR+vgalPM03wXRkpHpa/iLo5K5PaUCmsw4HlgR5hfp7jEiR0uLxj/
7SNfzryAVgDx3gRRgRVFgvAER1JJAprtBcuTGQAf5rXricJoHoLdFKq4NHZif4yz6FLt4l/oMgUr
tl/UgAv+QQHezgBIzVFYPt60b7zSnW90nbxbR/ZGdpJ3i5oh5fV3WFLOgt0Rxc/09Y8OiJ2FnBBX
ZNlbviatS/El2/A0I0pN13ial8Ye8A+vNaP5RJGZf3tnXv4QFJilc2SlCoxcTU9zguODWUcrI0Mm
06dWN4M55oLN6qSGJB/9N0Pyd6il36S0Tn9CHLdHKfvoSJ4M8ZJBy8QDHrh6u5QtYIpy6hbFZgNJ
q9WTBKE6oiaoLfkpCiNTtYVHRKQycqzyyc3im38BMKgJPv8/GJKKSmoInppj9++/Yn1l5VB+WPhy
8JIXFwq7G2TSwCV7BTzw/3OrndI+y+BgsMKC81iK1t/foJrtuI2yFCgIZ5V3H8YyQT67DtvLvjBD
ixt+bxAcPqNZmiCwiU8KpVr/wSCB9WoFI+kNcSgqWP20sxdXj3dXibOzFKpjOAhxfjMjYdfhWWA/
kCVSjFRPqeZZXQ9ux4YUc5uR6x6T7eseCPhftekszTQW9llSMrcYETDDV+6soSVXNRuc2/t3Yswu
geyzxq5KlwFfX3Wo6KjsMqgYBC9gMYs8SUGgT5xywv9SPEEtbgvxuYe8BMFAllBmEUA3eaoGUZdN
NVVHBFxKTO1tGCy0blpgwgP9tDw8gyVXlvHDMnwHyXhm4K9MsecxQwaWjsW67y7+GGkpWw6V6v1C
Fnj/xKw0gz2ceM4fNmvKPWRod6S9migkeZt+q7VX8e9nLm0HR6O2HsjbL9pOHIWaYji8m8Rr0DlN
3KT6kGcbWmqlyT2ZdZXydCxRRJIFTEtd2WJudqwkFmhATWVYIqv6OYO06jfCNEzGZ5/JCOffFV9B
RyseoGRQPiuVYb4CK+5J6shi/CF9q/5Q2hpx7K1ibXFZcvURws1Kz2A7L/h/jxleYLZUaln0YPkD
7f/a/F/EqrAzt269LjK0pRhUBm4jUe1eBrOeuPMBg5fi+ikn48vgDOaaxTjB1zKD4j794GGjzXei
ZMz/xSDTU/qcZeWJ8j4muheO5WHpx5u0mJOMOkCgPfsm3mIhd7hnxLRUSLuYjtl1mVm+bDikpy3g
gleZ6dmun0NuoN1YUxn7VjG7Cqo7FuHlzajKllYEBtVUjRNukaeQMwZI4gbtBY8AyZUbEw5PIGrP
9vkhxWEwPZW4SWXJE0zOf6MR6tO5DkJs7wWz6I0whkhDwLpmxn0yF9m+3LksWnty/uQGwKIU0Iym
gVLu8y35l1h1SK4Vb67gV4q+tPTO+1t37e8dumJ2gJ/cA6PUxzOs7vFJseh065mrK3EVDWp3pFzE
M78GZgZ0DoJiRicPkdrm2AA4Qlb/KnLn2HgiCV1olW6RIpM+JZmCOe5DKskZHugzVdSNJm2AxVBt
sZiaZqixR5hbI86+4ew/V4RLDv/4nDK46dBaBWT/+9kvo59++rZKDdiJQyYj28Hq/3JEJHiM5RMd
Gwgo0qFUZ43o82wdiSjTpnLeU2F/GDyc6W8k+679SOR4FxSkl29jBPZytE9VvXSdeLMUwr2PUGlz
U9BgaVZTRC6uG+klJcIfjI+xeaYTL55VEFr/8vSgXiGQTxyG9pxEpApX4dEgxVShRCLZhec7A80k
NVQcq3pafibTCOwcU3x+QpdYMuOtEx6CSoKJyezYaEffXDFvv5KbeRGwrj9w07kONVGTMl12yH5l
dBBMxeZH1HAmnB8IYw+BXI6jICILiv8T/dzmx25/ef4PrCtl+64+h+QBYRG8jGUBwSGHUzBz6PFj
+FBjfFmhlqF2PjAQrsxOLIWqtdiSV+eQbN2fsFU0ppaZr/XxhxaiEPJJ4vPjJcQXUS2SesPZMSYi
gNnlpsnqhlpnNTEpkVzVY98M0DbSWvQGq0qTuzw4p9dzwcAToaRBTsHRNgDZd8NldbD+cTAa+Fxh
FW8v/6ljfUwtV05JX+4sPfIMgzRqOgFQoxIBt0cVoSbpCK8sbfF0bugyrE9GAUF/8gC0UETh5dww
PAwLD5Plg3FzAXvGierJmHOQK3vSdG4otGW8hAzhIr84BAkS66VGmYZiNMgnjsQViti8+Rq3JwT+
cl4jtHpgWmk3MaUsFQquD3wBAtfi3I37d4qADwCneDQdoTjWTlk77aidLPMP9E8WFanljwLOwxUR
qFk1kmN+VSuJqDeazhLLVzNyb/J+fwHxB3Rix9rOiZJuu59sd0vCmPnoDwASPJ2nfbBkv1KAk3Bh
26kakleczBriNUOxp8ChdLcHRzUFn8WiNUtUP3pUWthvc/Be4WWDaZKOqXwkY2OdKW4jkWoI6jLe
XYkBHlor5pxApHyHUZ4QmNRxRyhpIhpVFSSINHREoqrUTOjt5TzrpHV6JYApvwCaOlO2FFX3OClw
tW5t8ALG+yCl0I4s/FVZMWNX1pNJAx+VjN7+ZXXVsMdh/5AZAWkk9hm2e7TdcjvXc1gEe/bRi7gn
UJyIGpx/MyTvrXvV2lzxIooT1tCpM9VwMcxUtXJ6JluO89DkMWTH+3nTeVR0y/dG+nWfBnn1GsWk
/LmLAFdFnku8MnQQVzurAcCy1nX2YVKZB3xo1b/Vsurdh8mWM9SVfrsgZSlQ0MoXKfe6h9k2I+5H
DW4tfiG19RNuxsU1M2HsaohyJ26fxkQ2CtcTD0UK5uw163qmV70Mo0Fiy69Wbd10H177v5sK/feN
+H4kPGBW+7AS/03ukRYAo2egQzrcp1XRSq11W9GduyVrNS4uZ0aMfLvAnExTLGjay86ZPA2Vnw6x
8TOFCAXIo3FQq9uDfBOyvA0BM9/z23CyFMTBdF6aB2XIZ7xfPpWSTzz1UWaIQ0o4opHGM5BSOvjZ
RADdzewwcKeR7dgo3WejKUsOXmCwvO8a1fNpbA1C5QJUdo3RlFxoq9EH9B2wl3KKKEjshDvBsA+9
UcOvdlb7tj5Wx9PPJZ+z2P9k8SXj0n83Zdynk9ezKTucQD5bhTdkYncyD7oiqwFifWXVxVbOYn8u
8zJnlh4NECG0jsv57lAdXJg8DSIDQDq8QUtNjHXZWGpIOom57iMLR+SanCX5BOzp/MP3jGL3D9Us
gASDRO7xzec7coYr9U8xHYDLODnkLYUfSiKJc53CjeSUIGUhftQtSc7T/QUD5pPXyOMpCPPwG8nv
2mVCt4xrbSrAPIV2JoUhbmwSlrLtbjnqQ5Vmiqm9+hnI0WxBwjcKAcWc/GOzWgRddfdiNBRorTlg
Q4wDo4SfXjjX9AUsiqjbdMYu7GhADA9WEwUrSKEl+biM2Z2VCDmneTfBBvmazSDBso6Mk5lmsOj6
CsNE/PVnN4HVfWj85mvRJS7altGhEiqfO8dhasCcaM6d4aXLJIEgKDwwpCPXTp6mJgJ2Q57LEc37
P3OPkGh46w7rE8a9K/5Izj8EbYIR7JVnYBqGmSdOGqImgglsiKO2skXKYlIiqhu9EI2zuSCXdMJs
Sb8EhqMcoozUah+CUwOrJ3s2di+YwpXIYsnB9UZ8UOafi4+QkbmLPYekbJ6wKv1eXdcQCRe9UiDG
zfX6DlYmEOzyF6dGu243r0rPauO5hNIr72Zj7i2BEWxirbL4Jbqslolk5pb0aoThMDNIp1VdLOuH
boZ2M0wGZAkYgswLrNFmWe0kdUg7vqwv9uHKlowLEEIEGPTD8vpAaVwnHDXUO2i7Y7VW/RdxW8KL
QsZgWa9RvYMJDrT7/wpy8Rsf/25ntC0xdMI0Hj6NFAMv+H8ashUdji1tNHBUdTH8+mRWZFwD0ITe
9/KFAQo5EGTJ+CK+FcwXGIEUb5hpk4FXK0xUnCiJE/GQb+yTtpwZgqMuTUil6uDHXNzjOw1UYrEj
cKyOkuZ7QzFzcg7Wg4LzM1GPwhPvltLaNcRksdJzASVJetC+0527qV6vakWmVqDT1E9eqKo3MvbP
20d1k35t6e/UKBi+kQg3QIa8dop6iWPS6M3OS7b4wJ2r1cB+FUAuv0i1e7hlGuSQR2h3/OsbbP0t
JpyPuHYHIZBxiMFZvySGbCvSvvHUFfPG6WIFYEIe5kw75lnwhNlOXUK6M8kGPihutuQadMCuyEwX
uOHbpjMUp0bwepDiaNkqAVq8Ljd28LiCDU6Lyace/pjLNPopi02SEg3tbfZWO5WKafSqq/dVMUYX
5O/UtbwpfGuHjZPoj7BmuNj+13oqjkrvBSvtX3rX9L/IBkbknp1umwwtQaRw/onu+RaSraGFxucK
OzEbz4O3OxvYxNB9j1LgZeZtox3rL1k7k4MNIKIHzaQfgCzdUM8UgzrmOvGfCRoXFPx0d+9kMv5o
szebKYlDkuU6w1QczSx98mjCB/dXpcyQp0okyZ9cwqxXRDZscHc6m4SmO+5BftBj1vqT3wldsUDL
OL/RODgqx/Qt4nm8MBVAdJnVJ5sAovHkMoEZqF60lPUlrkeFrnqCfIFNciVT8NTnSljgfA+mONdl
uPL2bOXpt5as+1tUl+Mkoj7pw4qM976t4UPogilPQZjol0vITNs/QwrHJBFRiGG5cGd7rRkNrxun
Dt+weqTBMbyxP1zd1UWyn/J5sa8TSn17x/5t/76IzixpDJxs/cl9UTVnfVz4CH6u90MaKmCm0vQo
YdBlN7wunWVoyJjMpEP9zC0DrAOdlk7dNzF6AqdpiPEVQvEn/3zAEojwWLNL6uLySHEyjKpU/5Te
L7xYBHL6zNEOVt9nN5EESdQhJPgfqcK678fowxoseELZUWyLwHtDc0sS7RCpNf4eCrgxJOG7Tyl3
LqbfAKLA85gHDOevPiXXb17OWlx2LwbLVh1+0+KZbjLr9YqAdeFL8NeRSR33IPYI9xC8jK9faroR
/7xcHHlSubyw408j7NvrtpDYmRp3UaBdPpm0I6BloXfko/T8peoMps4mXFR/vtPrka77yAmSubTe
74OfVUkZo3htB3fnxAqoUAkAFHEPrXweOySDE26Q6npnLpxjKNHDNJCQLA+VF06Q2QdhWuV/MyUL
WVePOQttThEicyHitV0Veq+DdqFycwN3Fv5M3M1nIdTOIDGaub38PEblJ0DHByslMViq4ByOy+V5
eUgsGdvLz/dx55GHGefMA9g9073zRe551gbV6MTzYAKAkjc1AIB7zbPGNQqgmPekGbVsF1pu/5Z8
C23Hp1qvv30woxmRAWWYhnAeNXwdxExW8/Aj7S80sM50MXDWJbFxUYT5xJFb5QTp+bVVDSF+c6ah
Y/0uuc1mS1BzgYA3wbps/zMdUS4313j6lNixOYMctT24PDl4s3x6u3c6ZEGsflxj4cN4NPalIOTk
j6gedIU02KYJVS8HpqEVWebCraZ9KkzXH+NVNPcV0G1g0GElcbKcIY/083tMxXdJcHUGSV27r2Op
8Ns69bWoB8pPsKvAN42jxNgMZo2X4his+AsnqMgX0w80Qn9zuF6tKkamHmP0zRDCLJwQ/clku94s
RZ9OXWrIn2egKp/osXmoO2sjcXD9Bzwm10RvMJ7K6B4eLTrxnoSVdPnz9LDqWwRErBhVvSl4HA+E
aVsDdPsopFB2kYpNFjoYxN58yRid9CZCY1rp4lLZBnfCqJVTd/0k178fK/szSW7iJk+Nbtxh+3BG
7PF3vQZto7Tp3k9ZwcI/mgobKQgP24siTCpgFrn+Y5VSetEICXsNVZ/ZPlV/BZk1yDneA0A9/Wiw
tGyEEsJcCoEgPmMl2Fs70B4B/zresUzvvzk78D4q4owdI64jT8EMxQOmeEeLUznK7McFqLRRfXlG
QBGS3kjgnz6AGPHMdOA04DUlR4ncOBc5M6VapurzyqMthxB+SBsWkUp0CUrJzLPEao5hUpyPyDW9
rwjqGd/H2ZK5cuq2lZBdlPojZjw7LUxztyYAHchJkBEzYqx+t7Ygo6W1w1ybi7MN6LQRBX7ZAePG
BZ0kCFOZAMogsJ9y9gKMG/O5/b7hNyX2EEvIkKEbU6uotTO5tIzDO3zAKbzp03JxYZtI/Y7lJYl8
hPE6vr23Q9OWtwo3xlTWW33z+FkSdFbrmAARipjPJ7od/G+OxEg8Uv3ltpxW2YOqDdcN2A7lzw9o
POH/OH+khs1bdHpNKiXbwriUYF8qlv3fNjCkKbWKF7mGVUi1XQYx6ZAGBD0EcmrGtd1y6DCjjGPU
aIHhlcnMJ9r70vfGkpcio6yF9a9nBzzV27Kxs2Igvggox39x1pchZ+SKvrNZ0W7JZYbb9gpWkfw9
N5Wv+5dYHSmx+yUB5y5mh4JpJW8DZ1jpzXexbiAE5qTR6RARak0+m8v8j8E1CO/j3y2HAvc+evbx
7baNvY7X+iwTth9eXIYIXYSgE6phEf58m9W33OqVxYwxxt+A4tCUDckzcHcVZR06l8UXcYXRW3h/
63Nr4EOKKbjGKHO4k3ZmpVwZmY28cnJYXVTI3lsJzinVekYdH6NLLF2v/uvxvXWtHF1dzxtskw7w
S4XHdyDA/7S4CWrfPuWb0LPU+c7KKpYOXP8kzEbJOhCaKU5rflR7q5PjlVJCe1fufh0MVjQlMZvF
CMgdrxxlkBkp0hJp2KYoRBsUSds/HOuAOmjl7KibLyAtQun36bvKqOfwl4wA+tirs85JkZuBrTwx
pk5UlkMflAM3yic807qggzSau0FpI4f6iNGK/hJpcEYMV3SPtDH/rbxi/haN9ubuT/hf8jCSLREE
v8XT7VDXvdTS4RDgUyF8BdNpbDTuuPzk8lqoFAc169nJsYOZRqQLgdeGl3FYWqmGCmXPLKkh0Q8A
/7AivzlDcBGF3MKOwNRScase2UvFxCCD4EsFqxfhHR45JKhb4usDCaHjU/DT0CtUwcuDW37vMTcj
DlLhnD2garGNtcyJqxC33sfJ3/T8gUIk2RQtEaSaa1jVxPEyJfHcPvLSvMR6MfHaNyALmbGQEGiT
Ox0zVuFq7qKFAJksMOQ9B12ZxwnK0BbngcYa2kW6wvOAc23hxlSo+wvB2kemse+0QK7KhAkkhV7d
4FN2rLBWMXp3zvJFn/VNjUjuKHcUFwKJBs177043+gLnpN2qV8JVkhvB3ycCCZx9nwt+CJAKn2kH
THco5alIsbMInXoPfITtQpbKRSL5cHIOAHv2qcww7Em+0Gng0SFu7sxf/wBl8Ck00X53KMAXjfPp
CV4UJiVYistAyyggkhQZtTxwHVfxQOQm1Q5TlK/dnRgPwS4cr/Br4rzfwu+1a0aZ8n1y77saST1W
40I4bTs9VJ0AD/Lug8mLkgygZc+OPGkBhNehUGY8NS/CYlNxGXSnfGMjcdHifUPiqCcllXxDxrOe
CzG9sguo88ZPymd6jVcZj7/BuetaMMODNGDcYMvfHUG9KqajtE23dxsObEeYiCJu1GrZdTVn+D4V
19vDJrAaRnLRV6CHph2L48VP74ZkdWqZp+dhlAGKJ4SXBZ4uwlxAYgc2xS1i5wr/8hh4RlyElkBI
GvbV6Bra5SxBU8oAAvthu9acRjmWd7Uo7PFHXsbUtHHCdv2WRvXVPcAqskbx0m3rOmddNKjpgFo6
qbZtorJaJhAjGH7dtwRg6XZ4S8Rt2sCcjKJ0s5mMF/xihAKhDcgyUN3iH4K5bACy5/Mse3E2KQ1v
DgFd5zMkwx3/cIsfMfwEb6+9GHabH8qbwak6ALaRJoWKEx5Xu6RcZBhm6yozl4fQyiax7T6KwB4Q
/9OjpMmFSk+jNm1h/RVuV+QG31lGbdGNOqRlkZMXWt4DgmYcw8Rkzls00FbHriyoT4Z5QnZVMPH+
NwPiNKEh2nI34IfplHfjShb+W3oTsjAjuEGJb6S9elos1pE24rP2kkj5PTiLHs6wwwcTLU2DMzhB
Ebpgy4pNrEMO5t53FRmK3XqO0k9So/lzS59ONzaL8sCqeXyU2QqTIRRa8m9p9SpTyT+esSa3CHEp
EX/scYuL55rA3XQXswJ4O1fx9adTlINqG4ax+V9gu4u9flyd1wu6MCr7amYZV+M0Pn035ELyfnzW
vGe5ErS84IPY7uM0XAELBIaEp6I8csGLLMlBs/m5KD9XV192m1wESCdSsFh8lP+QLgbunsmpoiQy
zA8Ypjjdvlf9NbVBZMCDrra733KYdXvr8pnA3lVc5RLzvcMelBhAfQL1s3JiQtqq45wCXh0i1J8D
4fR8D0hbZT8lxclaCeR58IfQ0rUMXAH6y3Eq5Zz0NgZkBwmmJ0w9CPrZ90y2hX/ioDF6sykpet1A
IxvEi26dKH514pBLCy8fBqiYH841UuBmoaC+FgTYC7g84pIAbE84gByXzguCzir4ip33wCUtvLiM
I2coj+Ge1znCC6WFFEu7c07xq6xibPKBPetmsCp5iTd9nrG924pFDrR9vDwqfIROwbeZ5FUkj4pr
dJIS9MccB63+fADJimLOaJzR6+ZwxD9Xj0O0Qf4kEF/zoc6wSZuiwtzgQFyB2vesMsmoqTnwaPvb
5SVBjl1TOca+XkMKcSMXHTOUCxd5/dNA5D/CM5PfUZ+gElUTOLeHmjHLhSjnyXnicWM9pS/J4cEW
+95na6zkT1lYR+Hpsi0WqiOSSknkJ4nIXKxGJZn+PARzkNoww+nV44Q1o1iEvmzcEbUeOi0LePU6
ZxL2jstGlSh+b2ZsZgw/A1A8Q+UdPaZD0KWYWDPv4J7OCc7qBP0WV5P3zlX+22SHD5zYFlVHUcTp
8a1SfxSm0hYtFE7VM+lDtqnjLgRvhuKVyZyzdRT5gd8VMAUgCiKoU4o4v8itl3sVbwOJSKSF1iHf
Vqhto+TuHUZ/jWrKTnudTM5jnO209fN4R4jCCa5s3C/Uzl5Fcef/AMv92fBCxwEuxbDIP4ivr0If
qD4YBg1YyqZ8ERyW+oZZ/uR3mcmOJBvmd8YcKLMVJrcPj6uih9ese+6fG24zlUa2mDhXiCIynezS
S/mIhO0fyH/RSEweMMTyyFmE1xn64OUT1a7MvbnAAEZGSayQx0uNJY4vwR3NAiaZ4BF70DIu1i+2
pq6My3YrhFp12AxE7t6f7b9ghAfcN7jSgLjP4P5srtF9Hr4pp2XkadvOuA46d2p0K/X4RF9RJcr9
xTHc8vPRvtyJ1/vqV3vLXNgnbUUyqqJK23d3m3hgv0FosGhbg6GdYRqj9d8XgDddF9wCy7WiN/7L
ojnptFjNDFr5ybF8iN6olZGP7NT0P++4osCV76OSO8wb3QhfXREq7qRsBt86gfCZmLk3bDaM1Aqs
2aRg4AYLTf97NmFTo9e0zTo3HR4CfFhbaDYFUqw9zFRELzQNd2dwhPROm50CcN7lv0uffITUCxPz
HVT8/hmw9hfVW2jFzioYpE/csTKxH1mbbka4pUkHVKZwuhFxv5EMGdtojUnR5lKXNUHQgRqinIzS
K3pFaHHZI/I0NQEvYrdXtjyyX3da9nLIPUVpNiUzJl+D5GbuEvsfpso1hHl3DAPRgDLWMHGXMghD
pOEXMipc3225puHh9MRWnrDoGvBztKM0rS6F5m/rtm2UT5guj9RSdc1XYPJ09Fug24SjFI/XykF7
wrX9MQgeIqgH/Cl+PZrS2zNJGIsd8KOYAX5U9u/0o17ia05/mVagTLtnaPycjKYaCh0Xj4RIGikO
VaqxDgKPCifDTaETXkcRMJO85lqO6aES4ScB/vpsruA7+LrBuxn+Ogt20aLpVWliv9PcFqtU+BNT
XR/N54/LQjmf809L6T0UQWMduaogFrkmtzBB3WqH22driI30oxTOVSzEeqc+7f8w2RV4zP8v8RT/
Z7kOXr1iHTlxCr+9YqyXn7F1Iw6BQwi2OYp2y6/m1lU51CaFIIKLq5i28BCdBlt54Smd6uxYnMZX
1BnaPQnA+xa3DjJzKCZf3NDNabteStJrFm1l7cUU4qkraLqQ+vqK+eCPs/zDrJ3hlh7SgXhFTQmL
SxmJa7jCK47ant+IUV7QyGCKufsoizNdbjeM785PrKklzgp+hV4VSJdVylF8m/IJIH1vtvyUZoDk
6UwbImxI78dyvSdqsVb5mXLdbBlnyWLBIGecp3zaAseioRWwDwGxa165oJGXJDOFRbP0FMpu+073
3YY4ZKG9kKHlAApANkn3rxDDSlgzgnP7fpAA3RrPlC/7rDw/CkMJc8xQFG9XGCHak2wNGXzBC7xm
zolCoYKddj7vfHr/7jBHQerp7d/zEDkzKtqyuFbpDAPz+ONnI1gRdkWqwdxE7ul/yclcdLqNDHc6
oafd9943dN541Mvnk9XD3yZ4iL0XiD0HiCuJn14pjVVLirEVzw43vr1bU2as71EldInRf+M1y9sJ
s0DfWSe2f0uZT3pIa19t0pqxSPFlVfvEBX6HV0YaEJYH0hectINoQpBVYZRwlWLVQm5zfcqWOPkY
GPa7NmIMJC6b+IDTz9Yo9TKQZveBRmpoopcOCDiZVxIHlzuIUrYunKNP3d91nlNhKl2YQNglRTFp
GPRu2Bw1b6l+YDtvb3mcXRLLtpLGQzzaATWLoXqgwUiOA7CFA4WOamcYvHoXOgat8LpxHkmhTwqn
RDdgOq9hiXld2p/eo+v8Oq4rH2X+L3K9xK7NP9Fn/lwDRFD5u7QPanWPzPiRlpexYBrwl4LXwKAD
D0+E6W8y+u1orKfGbEGmuS4Z42CuXgYk/fT1RUV09ZQsF9Z12OsyAN1e+PSja6VXiwF0dthorxZV
RnU9meLtMcUgay+KGJzeDFErgb+eG93vpiEGY4S8HE3p0hEm1O+MjiM94SI3Mv2wCRbW35ltsnCi
HvBOgSVih2gdh9Rwp+2rNXTSqUhL5zkconnghNrsOyQCj6pWLd+fAqQ1QJl5e8CWM58gO6iATP58
nd45a7EY24w7m2YsYmypRWuNQRovJvioJ5Hxnqg4L6bSnqpkktmuoQKiIeqJuYtPBfrxxQGPUR1J
awWRhzetWHFKbSTrLj93Gsoi8HpAg/sT7gcMp/W9sJFcQWFd4nkwae0e6y7AtR/eZ4cCA5j/vagO
BcUhh/NmvQIdtDk0akPhjZzsBV4BbjTZMGQBjGiTIg5r4vmrfcLSrqO5ATzyu5lLIwsVGTA9SCSf
HJGMLHtJucq/dDxVXU0525juFk40LD9u4Ygfrhvre4o4/uqTY+tuHzIvpu+aXHetFCZ28IFf5YeI
I+Od+4PYZkuVqSe3/wHUpRp6YSEddP1g1BCnHvUs6/BXmprRT+qRjGmiznKPNT2PajAZb/5U1fce
aJoX0UQTcaLVllLzFnCQSqaeD7Evj1ZWFOW5OUedLbxLivVQ/lE1ALlDZXNReMfxi6RlHR72hDkM
Lo8g+0TNXsBXv3UHz0f2C54BAvNPkzSkgxdpypAp54+NuPXhuJGYW8SFhAS1YBLntCgrSC8H21Yw
K3P9r2VUvRmrEamWs3ER3o+CL+dpLd+T9QXKuppn1jUHhqok5AXpWmG6MDboUALTORWoJdVqMWib
ge8bonnVd5mFSZEWQERGjdyQnAvZiHpgnc2FDzjmggf1P5JcTRFZPwUQsmWagFt63183TxoFzkQe
AelTWRSu7qvPf4gWWN1GcQ/pAh12JjnRcxDEqMS8CrdUHNU79ABvM/7xN1P2HV+kPAt9aT3w3wwP
BRggMhk5rp591vBpbkLdiCD4WWl6+0VEC+KkWa1SSpupdLuJzKWHowMLQ7VZKR/WVIX0wbfDVlQm
x5Fl+7bsE7SeE03QcSJ5Yw9SkdN2ulGu6l6Qr/tfjjUpzc6QX1JiJj4qUjaGs2A/582NISKV9v+l
OHTPoRKnT/zqKwglmaD9YIiHOQJRu7gBPQTR3lIj+tp9Ze8ScSZ2ZztMQEi0nNc2GJ7501T5YSvI
hnYW2+qQwEsqj3y7RbM+reK1RqkuimCxBiW89PkfbA+SgLuJiTE1f71ib58Xl5g8o+eLEm5y/Rsf
Ut+tCR4TNP0/14RhtDomjQrIyskpSqS0ZLNVLC0Q8tErBFgLrSfTKF+ciP1QD9c0N+XQe326YZXj
gPK8vN8xlAGFWDAUPPJ8PSKNI1IWd17ZmSzkHyY/a523qdw1ZYLM153VG1QELeExW5rakICBt+LG
XHG7IZ6VCiFAQQGC6Q6V9jAiAi+o6ULnh/5F5UdJqrGwttMqGnJMUvBTW/MFyCnIQ0cUF6Ounylg
nW1zpaIKTYTjmfdDz6f6OHMD4PndaZdgpSVQptRUuFTFxb8QO+UAK8BvPpoBfoEsGP4JXMv4sETB
Jo36Sbehw7u+QXkP9ClWhhPJMYrSk8jlDar1fUbge8aSG/bV+LY2vha4s0BY5v7S9mFf3OoG4JQs
UYzGBBXH1fKurYRDeZFFbTL2h/GxFu2Zf8qxBr37RKtnGexYbvbnlAH1ffrxo5cSWuCJnXLVOmZ1
cvjjvWRA8y8FnpLh9aLEdJn7al4vauwMwmPIlB9fM8/7UC7oqWGTl5CQt5FHpsK0J0Ym4FLR7CKO
NF/vpdcXu7lmM47bs94z1hzHMh3ApZJ8hXtm1zM2hXN3hxx7CIv4iuzxAp9Ij1qX6yl+pd5SFdwK
oBnYdIaQMscF6v4vY1fL7/xZiPYX/Usxk6z6xHo2K9QqK5vdq9eM93mWy65OMtyfgQddF2i8Tf1F
uD5erZR9nKpUybsy+X6PTL5m7WH+PHid2bw17AzwTin/1KIw+xim3wcjnJ/nR8YK7QKPbCxQUghM
4ro2GOhoFINR4iD9lpD9h41hIHYeCkS0MF63YUkQsRFas0bqTcDr2oe66NJK90ui3SJpLwrpJCdY
4r88qPNXQnUwA5i4tFbjzO4mcIqHCmnJXRkHVpvzZU3PPJAe5OgVSVBHs9ySrTN9+DjlxXXDaKVv
veDYsWYslVWr83YSfW+bWEOlHGawQjf2pB2UOTQtyyqS4IQhUVZ+yJc67TKJoT5jAKVvU7M/pL2o
33segat9XP8P9S/vJ0OX7bCfP8SXic/rWSV1BQyJiEHL6qQI+H2MODcDg5no5wmg2mHOj7w0IEYr
tKO5/lGjP0B3Y3dpE8gg3Wpp9OyYhPfWdsUVSSmkVANs87SsHV/dPmWjfRycEdmeU+m6ggevY98f
hDRkLiHOusCP30yhTICSgmC9RJGBZwZUfnItwrTrHRjMRR9Hh9fbrXUYUbVy1Fl+u3DCa2U8gzq8
F4dx8szHeGbST6ZeNELHpGWXJJ4DVOYBV4O8QN27njF/c2Z/WP+W2vawLyVFtwAKUhZSApJubHU8
lfBCP1t+5sDKW+ltTLxZfEtJozbKSf2U/JawZn52tyVTnhKC2a5fCOKokM5aktMbSmMLTc2F341E
/5GwjyRLIfaEfKs04a07v0Z+qWSIH/0i5bmXSe/ymAGx9oaNP+9bDLhXqEPZZqvLQNat5MHUfBBy
e62DFvNRZHd8soHxcFNv6noMeX/103ia4aP37hlTMKz4c8J/Y6JyH768hfHOxFFeulmq8bX5tVM/
hVXKzwYzWL11epsb76neZunSHjY0W9J8wnWMY7W9DcFdMrVRWzMHa/PwrUn5herc4AMTSPEnGDk6
fgXcMH0kWS8eV7NZLL/m8R+ai8bbePoagC7LruslNyaa5JnnypeBs4J6YtpULmJsatubfqJXPpuo
0WgF6pJo6cJYkz+sRHj5oEhfApm9nY+49ZBJwDg+BIyl9h2lIQhBBs2BIOhuR2XrS/GTUbwyLSdW
mbDykDKBuDDmyfPT/PIP18PjgBwdgrvoC5VnGfsR6Oojy/hhLhftUM1hwqZD49eat1MFfhK45XaM
r4o8VlkRbVNmvOiZ9uMuag+Vb3H/F2kbHcoTqby/gBk0Op2OlD9komzRL3C+YjqtUhsNzS3UIsdU
WHhRfrLk2kT0xoSPz3svNkP2lOOHDNafMfbF4nYjXUeNHowiSt+fDPhfgMAImbqjyYB8XLxxqIFm
RlGqDGPNAf2z2xbvBWXsE1XN3epJjaZGaO+zkies9ZsemTJyRCibEKoqPSf1CQWtGylVhQ7Cf9wN
IMVcMaf9V35aJDCiiSSG8Qi/a1hZiA9DfUKukAscDivYEXGEhjIOCGXPIOS6zYQpD1gmH0nAMOWS
2YLPZswcDqvZWq3vK/LGSo2B6osk+jzHawBFBkfjEE1mSyMkCMzp85jeOgLRdyocPGURpRKkU4mp
6yt2S7YZ8YmoAa5iKCm30Rcl4/WqeFl6rLU60lMuBxC5sLDT+Q+IL0xrQKqrM8wa0mr13ELIPv7S
9HmuZueyuk/ZUA8dG290xe1m9USntxj3oN7kgnXt89ydVrv/PeaAQQS7ai8IcTNcbtGuJxegO39R
AFxHrYSY9zfq8O5Lgz2yJi21dIW9v1ijpRaza+HZjYs0NvdQccue3C69VjZuJRduNM3FYUU4e9Zw
C2p/nRQnZdxm/wYHnJrE1i3R2Tmz5i0TrfTNLlmewXNHWwGIEPFaNwpzAUeFN/U0l8QTbdUqdoke
d/FvB3sY1wurpydITBB5YHJeKqL6+wI6BAewQg+PQBZI86yIA0ugOwt5W83T/jVMRjjzNqz5BTDP
ZiokyAPWJfzcayzWhl0XAXiSZm5c+KL7EUMil1aOW+vXgiEcHoTp9NNbz8wRpmB20bjXmPZ2B4XR
A/Pb7L5rAlhnxgQo/gDM3qc/PV8uhcN7gsRk0FKmRTa87h5z5o1bQrAdRb/3lUYM8tYP26W4Vw89
Lmc/r6DnvwK98PGPX4zE+h8VGcxPXuf8MZ4cPwnUHTsP/ouWJ16klV5hZldZg560j1RRDX72j+MK
ysTDE9oDI8acmhgRcEiE7FVA74zBcCQo9JIdKy6/qqXBsUH6tAwBglphZB84X7mcThYUspWgDdbj
w3Nk8EETUS/zjpDVJTapr45CIvkKcRQv2PfYw0ZiYdyD7NIuwsAUUuiN5C9M5LUZmLYuMBqTxlFD
SSD/PCeoe6Xv0vb/hd6tcZfsVlTOplA0hHV1aonvJ6W1onCJP+jv/e17EK+lJA4XWlga6hW3bnSD
U3b6DJ68GEttEucxH93P188+ZzP24/DmaANcFC016UvA37yzzEziJjSNsLzMLkNpD33l8XvpWZIq
o6NlrAmv9/703Cw6qOvaS8tf6xhjgFViZKqkgEj+/VhiPVwezVeAwq81oYwnUopFHPwmATKoIrD2
N80eaT90FJND5YnI5bKTrV9CcDGcBbdynBUI7cquRm69QwZpHvJhJVz2OxDq8WY0wZQ/0ULPZcrQ
EMNCoEcZkYDsPFzrh3fGtmkPan5MBfjSZCCBcAMpaJ7S/mknD0R6tET4VZsxWHqPxi+TxWx4dktM
oXJWIun23I13D+2OInV4RYl69h3hrF0IsJ5h6nTEeK5FIMYJZI/X0GCxShd0/fLmpaDwy3spDp6Q
NvqURAiEqkyjggaqwQLESmjzXzsof0lgAISaw6uYnjZMzB2Nzv0VRwJ6Vmux+gL/7JoBqMGjZfLB
XcUTTD4iE4uQTR6yXJbHgVCNWZGfcZBI5Oc07WU2P2/6TFytzI4YgVei6ioLD7+7xqYDcGIg/tOV
KbLzJ9TaG/mwxUec65g1fJnFnVG5yOpLEK122R2psUmITfo+hYlkzDLtdJzF6ie74GBEDB5qKpMm
eNn0xHeEI8RuDPJYjXNcmQNShMqPnesLPBP60ZULSx9lsj44nrQ2s7AGH0nhtYvCLXB3Wwk1IjR8
jhMjzumCAl1+vQ2HpioeBS2vzftGfbQdm75uxKwuUEHFL+JFA8hsvWSpFLwvvfd6l4CtGPUlm23u
dzyvXxM0pdZDqbsFiXY85U5tA4NB7jyA8XUOrjoIn3ijato5UPQCu3Qw6R9bccYVkIV/vW0zFUAf
gkjAshRPeqJT8WGdLGq00e09Pw60X1TQUOZIm3UCxYvxT+Jf4Xht+d5lOZ6hMRrMwfBasVGo6jg6
qv7iVu5EZPErLqP9uisnl+AxYMFPJQ5G31Fwd4XXPtRoqCQebmLaO5IS04FgZj66B+6g4EL51RKn
039VDs7/3v79DowHC+VbZUrp+TRjMVYtVnzyu4S2FUXlcUDbecCRg1bZBw2PPryKDlB457JU7GXg
44JevSb8kpFZVmpKDUGtVRmzfwraWNWEOtzsNly1p+AIMm+0p4iUXYijM6ZnYbJL2ftHLC2wh+wi
A8jnzdVsk0/aiTO4LVbdqa/q6wuPncReE1PAJGbg8sWxjs0XlhXM1hk9XicyZiCwVPqQvHZxnsSN
ctD5sATuZgUuq81GCkb/s8jezkR/fUN3q+4SIx/RlMhYjKLyzy4DZvzhbFurHIsZ2pGtIqIqyb/m
f2FB8ILyozohekV8JQ4LpdCCUhglUhi0ZRAYD/cvSQVlKhyAHm/vQ+Io95eMTCj5OaqOHFSIc2Up
2TAgvZ+6fSr20uKUteXCb53VPnkoUaFBP31BGqQ9xf8JzitHcceGFZH0D4Q63FXKLFdvSuuMO2rp
HViCKCVQkykju7pmljL0e/tXFG1TvIP2/H0t2cOCnFg4A0K1tKYXrX+iNLJQJ66JNJmOuHjRZw4u
hA1uC8tdS59XDejBlwbq0KQlkC1u04OStH5pDd2grmYIdoGBtkC9enq0U4M6rhrTFmcToxXKFrKw
cvkY6BtuHGbV5Mam5aI2WfqlnwLmmj7yRAzNgf0yMIc+ufyJ1WnLhR731b1t1IL66GEtMMnHUQJW
1uZQXfn5sLXtQkhwkxaoqWf1Meh2H8JtbVRBbt/hocJNOuSNxEUo8K/cYQZvG4+010Sy1jAckS29
BsXn9CezPn7VPYaAUUaMJANgMG0z7LpUVz6DWZowOamYTGz68LfafGBGQrRumD/8bXkU9xSPkRMQ
v7PX34srDqDnx/mOSBkc0872wzGLjsMOaBa1oTnACYfPoxORE1RHL1V9WpH0dS/xMBqlYeh86E5q
p1AmNEYjglA2tYXSsh1vE7ILGV2GzypNTi7OhZJ4olA5xUqIDyZOYGVNER9Pc63KSW96VJITNTdO
RhWi6Pun4m99gHfnj+cuJ0ZKD12ct8AursoAUGcQa3ZaTWVsjM1NlvP5VugIBD3A09lLfuFKZe2J
TiQ7Gt+o6LkT3yLdjhAfO+eELqx3k5/4cJ2ZisSbJcfqKSoVYU/sftN3cm+QtdCGPIs1MK5LkGvB
zf3i0Mix1IiIKfXUIESGPA3Jg3HAbFvXD68OJA7i9CD50dQdFg97RefdYl7Mvqt1u8YIUc6CBQ5d
kKJ5zrTENteQPuDseIuc5Hw2E+MDlmyOjSEJRiLtwQTQMj4/uNz7oQyXxQ0GXzVCWatQY3IaWvE6
CYLZCrmLgTICfDtQE81cZgNPIfwwraKeDGVWIAqp8x/hYBTqX6iwXBhe1jG2W9T5UhB9IiE0aroB
8zZnX+xPl4vxJdbimUtDrI0FnfJZsuj4MrLaIhbRFoMOxsQbZExRp9gNsiz6IeTyvQ2WyHR8tFAL
pLHLzTicJlis9UclYkyC5JCCBACMjAhkStUeIiI2iK6bX9POjkM3TGkN4VTy+essJE4FoMd5+tRB
NkMLWjGke1XkJ5pCdPs5f6kpb4GVUiHTU5UKc0qdwkVm41IQoqbA2bRxGCaAZD3KZWUJruwRUBvR
zMiauNks7WcusgADA6MkoBvXszA3NB+mym2azHN9kqPdGgyiMSu2rlBqvByLBNDaf3RaKgejHvKU
xa2nr+WKoVjxkJS+eT2Ng2wsDjZiigS0T2DOdIWVqquRguRHMA3MBtNCltuyxgVwtsuNz+jJ6lgv
edCifhc3DrLEBFLlVE6Nivzr0ige55EaB9PtdN6v79hw+ku3NXtaXYQgvM6joAzf183ijYgXkoWF
1fitvNJnu/ZXtOQjy+LS5S5cL/n6+imOV8Bd8c+jZpaH3FJw0mVB/omIuN9kYuUf2+iZ1sBsm4q2
bb40kz174BgLG+doppXhKATH2TYsxQQ9KU4qADRFKV3LlPxpM2EjQbbJsNjAuqXJ+dCCaqxT0E+w
29b5ENl+mvGwZIShDpxoVmcogqmqTMz8rNfqdIUE/PZj3ZVc3ZsQpXj7vGz0pVA4Jtwd085tuL0k
cJC2kjNIGyUPpnGcwaMgW+4RjIhOHCp1T5cCAySc2LyZ4ruEVnr+/dHA/cIdAfs5oiknPInXEM0g
x7mMlBat+zJaJGzKJzjCkfpkqgsDFr/8uXP2C5QyzgnK4tOWJi0B7Z+sqyTtTdv3ae9Zb0MewkOU
DrVIki2f3S4LbtjJWbNu/C5Pkh9O1qGQ/q58TfwcCSPh/3BZ3a62jXZKgcL/PJ6SvKf3etlV+mqG
d3mYfBbtTjJp+CEOXMPokwuXZS/8Cb2Nm4qDCQi+Bi9D5ndLfmZPvvN70oPWaPiCPvIuR3xy23U1
nR5p00EDdcXH1v0Dz8edGheHmNslONUuhx6jFget/0/hQAFNF8AH57mcHnHMSaqO/l/nztRGf3wi
vyTea+vgzqXdKJUxfvZBZ7GMlVyGhRWW2zNjD2OLCknIHzdX3Pa3Z3b6+LDOfF7/uIkzvXShqk/b
EU7BUEsGZNpeaNvIEZGuvSvr3KxomEVA4fHu2WRFr7e5gGBsexYlE/u0KB+Z1bgDG9E6f0o5ivJF
llymFJyKq6PUwzONmZ8mV+B2rc0xHjbd3xcRqDSaTFnBwAVJc5i+8NACvbPApfHH30dL1tznJr7o
WcLE9jbZccA56yI+z4lJ27iaSEhXNyRCkRPObqxsC0uorsowUJDNfK/r4GQKbd8OaawJ2mKzjtwJ
GnW60DYmMcFyyoggj1U9e7sn8R7eeBylnVdbqmSaCTQXK9qp6Hh6v99/BryspuQ5nc1AEey+ssI1
ktoToUsha5gZULuwiW/thiOkidDOi4mUwAFJEazbnxdf8iBU8CIsN7ugn4Dcd8I/avlPFL3whztr
c5ij8xopQOME5/W53JIOQIZh9C85ftDAaBgZC0fXxx3rbFy/PxKCx3eL/tobMfCnUU3O3B3wMP4A
8/T/aDUsfZ0V0XllqeurcS06BBtPALnAPW5wk72NHg6VPPJHlo1Psrwi6J5sT678KBoaIAOA5t11
YXxegV1ylUbo2iERqV3EA8PeD6lt3nymAt9aEs+Ni4PKVzUBXozQ6fLE1MP+Yfy5/3HPdWBv8QLH
jIZWDQOKwpNxoLJbMo4YZcjikEqYwTBCYrq0x15n1bJ/XoCh0yGrStBX9XYBVlgTJVs+S9ZnFqnE
WEqZ7X2IQwTqdjjnNBuqtc+neFOHpl2LTevO3U+PkecRXkMUFkTmcTrVjGN9+WFJm/nuekjWIZKH
EzXCP3expmr5LRPB/kBvA47mSUMTwaUlNc3SRrJFJVG/A/pqKFhELy+svBJsCSNooy/6qw8ujnoQ
0Wf8wRPhc9SFYE0X2LL4I3qOrQlZtQ6vNJthjF/xE3kgnM3j74JirB+pFnTkPdVGzhYiXL4wAakz
ty+3Atxs4qT9+ppZYEWZVsvh0yW7ZjPN5Huume9w0Ahv6DEmyex1BrwFB46nx094DCDss6mTdRHc
GxqyHm33x5EcwME46cYhJIu2YeSO5CXzCXmRslpKcDOBZFuEwxb14FmtdS9zRi3o5fPo8VgfWYgz
g0Lw7rRFztJRky5iSYDiO3wbo4UBj9tsd07GKn230PLKL/Fj7AfKRCvZjskaGxa+lXBdDsziglCg
3kYGeMj9Cmvh62nQUNNIbdFFcJbC0pxqlBxsVWKV34GiUKZn6OYTqkaBkk96c1hTxITYGjpJ68s3
pk2iTBxHXr099l3p9wK8lEhnB7wKCAu8R/JDd2ARFeC2vXsnNVJWxSmhv3p1FQKoc5aQRTLMtT4c
MpU1Gqlc4hq9SjiL6mXM0y5lSICjpLhA8Z2dkMjnjXV4sHOHAzFBdmaLegBj4AEUpUZIyk2GkMGX
j/S3vwXJ3hi4QalGL0ih5IL/0l1gsTgavvpCuU5ti0YZPRKO5//WCD9KUg2GH3P5QiWpJefeXEyV
EoFint3DDj6DeUQQ/tVtAPwnLpopjmsstNhUXOdScsBvyWrh/o0gTS3RhWEjxsdWrUCiZpMfbtGp
gcFiDMxoUBXj6QuaJesTEuHuI6WvgbzhUPEutF5Mfyh/aq4VZlp9B5oRijv1ksS44FAbt6LAN1FA
+WLuf0tKP4JsuzyX4bqEGrGoP2ctN7s5wV50/jBOl82Z3SVADb+6g4awnnmFCECKDIlErs9Qsc6t
+JI/7wDRq9N3YzPACjE3FRLfa6gE7NFhkP5e6SA2TOTRy54SX98VNIWhsA9coEiIC1AE0HRpMTWw
DUZRZ19NT9d9ug3Wwqr+tkHkhwcSMUDQ2N4XBXfch3Y8l+TF+v9vNN1GLHGuwB68GA6w0k+442CF
VcclkSjL2iZeqShY37eu9/x9Tijz65PBlmvjd9JqM1CsThalFXfkkJQXXwAcpAK91EjRmnBHFp4A
KSrHzNV1KXpPtLggE0/TK6Ot+8R6FxL4sT8biwu2l+qdyVRQAJuo1U4wrGEhsFtLJLqWwY52c8FO
3+fFRQJeOlKLEihFjzDyR0iiNk2i3Is+cuY6Z3T3PHzBGEMZ7eMOAvL2Dw31iKDkr7ZRrh6yPrqx
+mBYsQjenAR/kEUdaQ4xOZCPZH8TFZu7lpB0DXP+yYEajibcGODGx46fyHUG55ytFga7n+uSv1wD
IEdWzhTqlHw3NWVWfduq5RQec7G21Tc/iCWeUm86VFX1/FmbdMI6GJ2/IBCN/dn9nlNArbiY6gne
SPYk5ZXpZEr//CdYr+fd5oPOmieiHcndkunG/B05Sf8f6oGKN3WGcxE70bRHcN5C6qkoiPk5y14r
TTGEPLrUKkMND9BBwtnvKSpTvcNYttnDA5UL7bbHoN4l3f5gm6pFGSMDqPP/jjrYpM05b26AMq6R
PvUtk17qMrQt3Efh0fdlQZeOuKdP7Cju3kHtps1Pu5imImiTjD+vGLWeEPDFOEGbu6v+qU+iqqW1
PjdpOfQmZsu0zCXxeI0+WczCwYxtCTWxjqtJ4zdLU9b3JmSZL0PDbZhRTkOfoNmt8GxHSgngkBRi
HDV4G4Vu8YZfTEbI9PCDi+XvSIbMeQF85Cq+c7v9EZCnse/gtyHPgU24HWtMuwEHRyGq2BDJ7VoI
jvAtXHQyek5AK+aogLd2Vf+JYXfdLVudKe4PqRU3WCeQhhuDnGSupvhB5ZjZRbqyx/NBACVOHyia
DJ4KxFlHJm5m8Ce2i5LJSn5W49ceqX/wjGF3kL0m6N2Tii864+T9InvwD2L6yN6pWOaaJzGRPGHu
1w7vPAXwOqHlTwbMCjVYWBHxoIGkueltmhzrSgZvbDKyVTLFIECuWVwO1KQscpSDQgngPbJIen5l
jjIbfamcxfkQjgax/9YUoJk7/LypekW5yK5kdAjI/G/TMSbjTBLbIGmlaAO3yT361L7CkVa86kyl
7y3+Qsla3ZnKNbJbi/P2ZsNkLc1QtRW/NbLWSVUvp4rh3Ai6Tz1cUr/FrYDMeNzGLXYebuwAPNrO
1k/8IEYKZgsGfhlI/0HcdUVMrhqJJKIouZ4cufOTeGCpx1a6Cbw5hr/KwFx5AV8CD7sl3pWusJQj
NE0AR/jJDTudS7QR+56U5s+CAB0TpV2JlYmbIEAGnCJ/iL14uLhlsQEuLtCjHT23lL11Bsft9IEI
gIay6DcUnZstHU5X1FkzRnf2QesQK87ON88c9N1iAJP8dd+hNHKZFy2DvW1cj15rHgdSXM99HPK1
NN8Nqofk5VxNqIPyIpyOcVwpBqAH2KSNrOcIpu02294LIgITd4jQ9E0l0UmQ0pLkoOAcBIIzctck
MuW+CrN8pssZSZvMi4ZrYVfXEtfAIMqMTx9WAKeObjmkqY7XkWa+vCflDWlUK4cH1YPEtb0vJYyr
64xv3Bbr4m8fuPnUnCHTHS3kSfpoVhJTqa21TDC1IQ9xSP2LlWHCyswEZHVwu68Ru9QF69yYpELj
HaM2x0jzkSTyCqdaM0zgEU0uGRCmNvfllAx90XXX8+OYGDDVyehYcdfmqPYR/UNggqZWWeKhUH/N
k3Foo8FIZWrFbzQuiNln2xI7TGx+0V04jdD1VK9B9jQc/PKu+ikDqjD8M7UR1ZjSCllEg57dZmqx
0Tr3vV/9AxRJ3S80hCZUlU3xOczVwTB7nPnRklqorkZ6N9Cv7YONIqSwRf4EIZ9DEFZuxBP4Gtxy
Rrwy0WHpzd62P8W8cTJZ4qz+MEiDJSxBzF0t4z2bfEak0VceOrJfFtPQe6xQzvkX4bCQIZ/yu4aQ
7O3d0z94QLfk34vSzTXWJQSAPrZGWNx0EsJ0JT3T9b2h8k1VTMSJHdGPZUaTpK6XrXw/mEDhZZrU
8ZEmAB+jCyFQ4v9qKIm8h2EVuStSVz6BBJ9IvVJa/Gxh/4MdtWgsmsc1BU6Byz4oJ66J5lsqlAib
j20HZap3d3WD0qxnIqaOve3KByLpmemxtomP+NPqJ/DCRFnVXFpCl2K6jUY+2tlvVgbxcNcxTO4/
LYYtnIPi17ohvv09VWxRYcF1rRmmI+z913Fhb3r2J103V5rKYC2iI1nImbC4zcoATUJmomTDRgyv
ijeTIUXD7NaA3ktzoTc/lUikq67GE8sbb6h3fSsdTpTBjw2jkt+R5u66yl2bYOVjCE3m+Hmrj3uc
JsreNQVD3VtQWKboNsvQt22Z6ulR3+MS+LljBcXoms8jr4ScD/XToHuuKm5pbyWemhZgkfuns6h+
lBEdzS0PD4zMKPoB7U2pdHFur3GaNAlHBY231kzZdAVxqg9c7fpfdxQZbpIEQC60sQhNCNCgNHww
lRcTRqLRgxIgd0ijC+uBBVYRqnVqGl0mImk3wAtyyZmbiZneY6U9osy9fSEhL/8/570NuAaR4Lyb
BU7Axvy4O1nLfOIoNfkOte6mihX8hq10155XuMjFSXkp4OrKkc4z4f19D3P6X2S0YanQDJ1KpJYn
hD5q+QvPZyJxaJ65GhGazoR/C+hRTYREi0nHB0RYpXe4w7UEUaCZ0lN9HeqJ1xWNdjW7I2/xKgec
r4Xxg8fsh51sAKO4/K6f9ItVl+WZZ3lBzPqf4hSDgxe+5z8HA1waSGcD3vcNO0DigN2XH9Cjncav
x/Xz0ZFx/rYdyIov0GuyiqRS6lgyUlBMzKt0xnpJknwozCdYsNQaDc/Reyk/NcyLcDF3Xbz9JiSZ
Tk8L0bmACk4oMLPcvmGtIaR0xlkRSHrK5EmCCr4oYGAm/11VXRLZopzOCvkS0pH4c1/xZAB4KBKf
8NyxsH5bMpuu0B6E/5+SVyfLzEZZmGainRIbF/Uw/ESBVatn2UfHPqeXMYtlWgb/vmoJ0BT2pzgx
48tKeW5MfEslux+eFrtc+N6qro6oFZbKzQnXYldzHVEtOycD6SUgHqg5TN2haeYdVZqByyTenhfD
/wdPbh3L8Om2UjSmE8eio+kRUCcJaBhO3t45YQd3okZj2lcLBOWAtJZ206b21hT24PweFxmycmfn
/oiPc9Qx/a2NJ85ZF3IYu1ARTmHClY3PoE6sJA2BnA3JYi6pzyDD4JPZE3vExs441E9b3FTFBsc+
wSCMl8EGYoaPcR/m/N3KCoG40wCNAy2Jioixbox25yxSBYIfhMZNjYdvCFppk1pcCN7UgXiSS2o6
rW8LQCA/iWymvQq0o0fANrMds/t3kGND79WUxaXjCKt1uJjXbh3Y7Lo9jhRcq1CpZPSRPYLYNPmt
CprC+jy3Iof1KBc/oO/dEyxmVdLvjsIyqS1SW1nR03uUTcYlVg1YioVjpiGkYCPALeju8CJzUjlL
t877nlyPKq6HmyEopho3N8PnzpbhGL2HOri4qC0mJVZDq+nPJqfToDoxB1Q/vL2sKS80OUEsFcJP
FBSR/tsn4h8a50fkv2myExgbVIkgybv0FkVFL8XYBhkL2OiMaOOlzNpsSyxsaEU6Zhds8L4fyNB9
QhdN9fKDA/GtgSv9CPU2MvdWJqp5OLvugbQyLegENE2PxLPB1JEtzuQ8MSy/SQ3NT3DQqkRUXwga
kC5sG6UdJKlOip6TalJanUrtKneNfxsHJOy+A3WeiYMM+GkgFm1fGmd6/sxogfg7+WAKdTJDfSo0
oxechhWxLWS9fRGlx1wt0opoE8WQ6cENVdaQ+ybqWKWbMdUMiKhihi41Q1USqAb3A4YQaWOFZPfZ
TvRM4x3QISlzAh52Wvth7UI6cOWwvRzQ4eLoRSNKH9Ll29JHEd8c9yPkXvq0MuZbCT21KnghedYu
4Vgy4yqUZjjj+7TXzFCOy+qu8SHjjn1WCAB37ewcF9BhNYsUkJeQ6PGabLswkwSomiuP0Yndf8m7
vvpUsqv8ZM/c+WLDOpYGSPmNMM7VdaWExc7wJ6styyrlhXCsq5oQRQH0M5tq3dvJrD3P93PXA2pO
PYDhkTnbShc1zU1ojDm2UB5liwlH9OsDgqzkic/8WfVLliwv3gsGxj1dP57slWKGYQUEXSHXrpzD
w2FaSYunFLsMHZpdOVJQLl8nlTJaYBDgJUMQLWOR84NF2hcTA5i/oixmC/4ZS5gAceWgZMVl+2zd
cURsBKsmp8LsreQc8OtQBME76VVXbpumlOjVUewKx1pGr3HYd3TaONuAzYNDhBd5ZZavvjlKpEGP
ItuMKGuG5O6KMtEsk4VC2pLzaQnRRLg+Pc3v8daARHeajLvKk1nbuR+94ve8hlcJW9Tn711apEo+
CfjlQjSO4TF8dKi60N2uENWl65LfdsWSPfQIm2Z3uDJlMYlNTFqLWcC+n0Hl7O7oBPnsByihrbui
WzVjLiwcuLM8qZ+PkSeAfrfa8bYUfbjFEXzWCstWJeOMNV6dU7tC8n3H7UP4MC4X7+QPsGEFpaT/
RSRwtLF3YJiqaTB5wWPWWKom/1/I1L0Ijc+JGSfhry78QdKOizBVDQZjn40ZEr447jrc2hm+zx6r
9SF8x8Oe+63vCzGOrCvAVeleu7q+H0edJZJTLVi8D4k3IN+4HN4L+nnKmFA0lah1KYOd9rwlsNjD
+SXfnZdPrhdob+4dGdttLG+o9eRz4rtyxwCyribV45fwJZSmCjeCMYobULf1GP3402uQWpCz39rs
/JnhU81dspfReh1Z62Cusl7nhg322NJNqQWD451JdgQvIDNvhami8otJnwc01pXULPQTLfZf8IRw
Ch/0rr/IKEgDffZH8SQsgjyC1sXGmXY/FZv+2nM72v2dwydOx8z4lcj6+6lEWOmbLvOdaKo1a0AP
9sCQp36UlYEf+9oCUR259PGzK0y6DP5EJIuyzwUQ4yYGljwxyVs2fEeqznyIPOY1uL8SJMcLOkhU
TapY+eSwa4Mrh2DGmqEK5iV5R/bYP6DRyojy/PBW9Pq5rK011JiXewHEbfs+S3Ob4W/HWj4zddHb
cegFNc9LxmWFrWZOa8AmMSee9127iI/SCNz6T7nr7LY4K7acRw7x7j2XydC2b4aZcH4lvimo0LYh
mcPD+N3G/EIC6mXC1yRCl5H/7lPH1U00s2ffQHpNRNk3/iRuaJaHRMei/5dG04+bDbGBt6AiTtyM
/acM/660bdFSR0ygfHAnmCWqKb0egSJpqQUuEmm3AacblGf93mhLwitDYMdaKy4UauNovWgI0KWf
CiPuN///AFa/eJFk3pd+ykWUe/gYbv4LFKfN9YzapkSqoAeI3lIFy3xAIOSWESvugCIFxomBMf5N
l4xG3RaxY9IA3Rpa0pMe6JgYoqK7yjvMT6HXw0g86xHAOhWmkI+UQ9oMwL9jCoGUpVAHsfJWSKxc
S4coTnNK44tT/MXhoNSvoFVq8Hchg5fCL5Y16+AbGP//bscKh+6X+1hITgSItvEDkE9dFTH1WyxS
54UeduDwKMGcqGJjtizVX5UNDzSTDaJUWwrLTSORd801IcPDPaJ7RfeHG8CIRro4jHGWYDMBCMs3
apLXkvVu0eE6ddbb4cvMoMl9GkgYUN5JozReKA8uspH+fJvvkP9ulg6pwgBUXdZbN7g1oi21ie6P
D1QuohQwOSoq/wEVQINJXTdZSRpq299+Dw9Qwn51d0AJooMzRx0lKpO9T2OqJ024IEOZ66gO22AB
ONlFYDyCPGfqmyaABaB1YYNXZE5etfADG+Ph3nufJJDR+4qd3AfA1ZTQ8ZollK1P01a2ieTQXTtT
VY60UhMU3DIpLdJEk5nE6ZNe3ZkhVmk8/rfFXvqG10UCC1gUJZ/zj+Y1jnuOswiwtIO0hmRr1Jdz
K3O1CKngM3gdlipj5hn4a8yY8hVixZqv2etT92L5eg41PHV+eBljCzjLp/V7LAk3OJDm6KAnkkzS
dugZqIELa+v7hcIGlDXI+mQHNZdrWenbgZqJExlPMSdBSqcf3jYI80XXIYNZa7GtGsWRnfPGHkkZ
+NMJHdpDHdNwja+4MSZqxP1pL+NJsxzZnIeatP3fO/q6uCCf7cJiNh7o/d0vvRb7lYpFL73QPpqt
4GrnitMX8NnWtTPF658nBs2+piyR+t0oB/1djtGmyiBH5B+JD971vPuKBkfkIHFePjN4woLB4Z4Z
UNLGh3rNRjdBXSrWyMlvg0G7O1+BEMiodoX7d+ZTALxaICc7fXwZEyTAkyDB7DTCMmu1XUK5ssPs
Qo5phB2eo4M/iyHh9y4ORm8jvFTFbOIbca4zKY6LcRI9u/jCoGJWUHgzk6P3+YM8qNpKofj8y0fO
pEoMR4j+n/QsLyFQpeIbwc2u+6TTDe4d2beFAN5PDqIfJzlqCH4EHQvTRMyDYgWIUTY9MG5r1PL6
4XLFMEuuDQ4GEgQblIXjmdU1C3iLE63JUYJbPLYUQxWKBOthFVvkaR7+rE5WPQ802MX5g/YAW6bn
UEl72M02rjNYYLlcpl6yV2fWKmieUFvC4giAt/TftjxU8Nrz1ql8hUMzwPhxlMxoD+IJ9CJQx4aE
1Tk2uIV/BINfqZRjasxs2QyXmqe34AQDOxxwqSv4p+aanFlBB04HdBntAImJFcZROTi3BaQCtR3h
a1nilfzX7hg8JkRrJDmHHyk5XkjBS8m1xKDfZehtt2MDIe/Bdp7UJwOZ8Ry+m/xq33NlGLr/WKfE
nVAO2oBqjSyAd80BTPdhZfTlvgf28GqhV2ParkmrB0OmPCoE1lM3xmRuNFzz6Csmrh4EACoTPDgl
uCkuH4g+Z8KuI7G6L3DivcFPTPes2qt3rGVGpL0YQtGjq5PZu87q41thjo0RV2j4xoXPxe5x0n5w
ETtobFJPnzGuCfpcgmrwV3FkNFAjQ7aTugmlixH8o8wCyyBZ2NuEJtluiIQg8eO9P5e4liEW0iK9
oaJLP5CKBgFSAEAjErStECet3H1uOLJiRpd19YozcIR4Hj1D50CgNgt9fXGKW422QsQoH42sppOu
+SJesuB3fs3KsleIt9xXJVIt4qeHMMOxyl7Z6Z8m55id+GZPmvnlgtAItV6fFOfZe5pNsL/1Ba9D
rAIOUJlk1fx/FQZ64Wvnv5tBuIoGtWLE+8GP21978bHBYiSK7+nUxevD+dvCfJWTnojKRyzbwdYG
xCljMX06SplQr7Vc0DoFokJEAhkXH7Ab8fotYcxZBcZEb/bG56Z0fixDXnwAilcNVjL2jCh3iXwc
Wxagb76ZPt1z1XKi0BHwXyFKBB72gL+U36s47Bd/bEjg9SVgiJ0ClAYgUotOpPjDIRdPXRQnLO8x
B+lL3F78ZXAUXO/LRyAH2Q5tvjXYzf9Vd00wHAqyBh1i8ouo5kJ5Oe4lx16UOOoAeWffryzxiVzE
7L0M898yub1HGJcWrJwUXYzExNDHnZw53/VZU45FlBgdAP5AdWOyAzLFc1U0wkSpE643LMxLJDYl
CQ2S06GymYhtzKDTrW2hm8bNpFxaL4iyL0ID9aKYiTUHXJ3PImFfaZu36QfVrjPRI6cvsWLO2j0N
LYWJGEt80fEkzgM0zK9vFeN+7FmOKv9fExrwZBICMXU6wVUJCv8wFduC9CRymsvICWb/69BMOnl2
1UWTzzboPvrCzPUvaEFSczS43oKsld16meVBQ7cYP41/PVp1s21WAZ8bcku2U5toG9Hv7s4jTBks
qz+zQ80RuBcoVbjf0GZwt/76m4ufUPfeeynelxSIX756sJ4x3fOUOkSwy9NoKJSBjjgAyFr4qNt6
K2KvHwnIEr+SZMJ8jBcOU0iEHwh4hDR9Xk7+wjxa3z2qUXdZfy7yYyadjME+vK0cZUCoUalydmxS
ppIqQCAc4kxvNdTJ1XlZ2XRaRGfwq0CX8Dh4Cd8xBAP1rEVkDYVoLyqryrONLq2nhT9v5kqXhqAp
KMRRStUYvACkJ1tZVYa2S/hY5Kfxm1EBtT5aL0OPIjeB/ayVSQdjQwvMm33BxXgpLwoIOWwtInIY
Ia7fvXgUKfm/nfa0ymSdKJ5oZ4rXDwOtNPBYAc7zE8I2KAAUyevzzNSYtnEWo1WCkE3U9VpZ5eUw
EBGxliNcyBkQ554C/xfQFWDQfbtP6uRR6WKpEGbClmG6c6wURFVW/5Cei0hjWiBdDcxFZri8Dpqk
xIPlR7L9MV8MGn14soCQijRRBrPWT7OWWZ0R3Csk8+HgFOS05XCmfO0er3lsVTU6AasKLeB4U6w1
YdTINFThr2cq95QsPQmDvjkoL4XYpG8HklN5d1E+gNcjhJmWYk90vb6KUSvLHHBZ8lW/meELaTqh
ns33Z5sV/h66mAmaU/ovT9lYoColkXedzPoC06tgFoOrT5f1QHhXGXzJA0qOSpNjiRl6ClWSkSKw
3cbU2eoFXD7zMY53E2Jjxr3Zb4mpb9Mm0kKHr/9Nr2r9WyJufFX0/WlJE+Ujn3qeWloA16Q3I+r+
NlivWCp+tFRnDF3YsBtah01ikEsaEK9bElJpXHDj5UHdvsxiWN1y32p0jD8CE0ubSS0MKrbMpfVP
G2LaJnTJMGVwc002aiLvzq1VwW7s/7F8mDJJOEpWcpm3I56sV+5iOfegPlXUqOYbKOrz5kHpnV0h
PKoQnuQv2RcyCrPgSzJ+EsqbUMFp7NonCwCMjbvyQ0uVEMoAWc8eIeu8vLYrnQQKNBXqVJl+ZP1j
mJSIAhJ05ppVJLIsh8VP8sY779rQsmjO5DGpDUgziPQ278esPjLlInRR6Od5aNZITw2BmYz2iP//
S14HIROZ8MjJgcaCTJIfttNIxnTJXRMHoGWmYjW9UTIqaQtUv7XgoD8yhHPdx+eRdwSRAS4OTZLt
7OfUaWafmESqg8tvmP4B7+2x16kAoq9PDafEBfzORpF1fG7PDMVcrgLqxSZndF840ppdK+EQ3z2j
6W0lZQdUD+8gmnbDZEQLzotFjb/520Ywz2+RvzbUABVMf0gR2p/EHwKYhEgU8+FEq97yPXW0x4W9
QVu6JIlSAiaqpAXE9y+BHt9JEpzIqPHDKze3enw0IrAMudbw0pcJmn4pc+2dWrQ5ndsPbj+kEZdR
CxEGS/v2pD4XCuKxAPZLsO+NfYckNcqUAJSsx7OkZucMbqiTSHvrLkBmMHTxUjy1jBmEMgQSzZlj
Q5nlWMqE+h1e6QzqDXqFhFD9bTEbe9ELNcDT5Jr5atYx9+2pRO8fQHY/USg0WkdW0jYDP78qLEZl
tC09o5wDyPn+sUfM1vB1RRjPn1mozcYBHuxBV0HajdoYzxJJVeldMgI/piRzmPWROWsWp0PBOYOe
tR1OuylmgqBYXoKmRlP5YWOmF2M9anXDVCqZWBSmUSls5mJTiehlHul+B80RNJhujuSDSftK3nF7
6wVFVu/k6He01laTp9Dj8gQfmICv/yzuC7Zy3+QmJ6GqeQn+TBQ/gwWHl7XzZq6QCwARkH/uV+S8
mCCpO7j26UKWFOXnuiuz3BfOf+UPrw8w9rYi3lMHMPAg3fD5ylQLiErF1BwM/edtvOm4ovV2xipD
to9MTVa9CDOMWaZdGVSL6hD6nRl+U8qCBikkLHnR2bjlzEUq6QlQ5xE0NgVkMej6eYyaZ9WqQqbi
wia+nHwa4Yz3ww6UdrGaTR1A1K2A4Tf00O2eVTcf/9gpwfF/q0C9O+PkEnK/Cgcij5aucz4xuNvJ
BeeWGJkM2tYFpbxzoww+n18jEGTostGTBmWwc9wkH9PskdBSLBvvCnT3Flv+IVlUB/gtWlm6cpuB
ynysNOra9e77kzX6xFkEoIxjP36ySUY+L918aItZ6uDj73B1XvYJJ2I7N/7g8Of2TB7lzPzeOmAU
duMKmLWlGgxHpUFeHJYkDKLtRlZx8rOVxCH1I6Ky28Bjk/8ld2ezuITt58Is1t9Yq6DkUmB+G9lh
V18yZY4yBm/X2Ic8F5OjM5O3TbvLvQRa9RSsTdIapLzae84gUxmwUfmgfGvht58pV7fvffGUQ7OQ
D105j6vig0REeG2VZOBERqlQM7IQz/Hmy6poWWZgw3fIUIjoOc/OhTX8221VTRGf2NuGeys3RQ7h
sdy0tPxT23LvATtuYqWb5jpauDO6K+0LJSt/8F9/CzPeMxu6T4Tmpv7RcZDdrwDcD0jMdOFjGWqa
zDDA3Lzn22DLeSgYbR0XBkbEf6EQ4fqkYAjw98bgwngyz87ZfdG1zSQs8Y857NuJVNkwlighs66G
dmGnLvzzvrHCGFHMMJwTBY4FmE9Wtk7DYMYYHEKlaXknmhyc0CVYViINusIwPZ2wNEAL8VdxP1Ml
tw6QivbfQtwrgZ8OHl48rDWKSCRztavKQi9k8TVLZ4FpUbctnx3JOR4AlzR8uNo7P8ULJAIIXlI5
3V9TX2b5Z2r8UsOk5ZGp35+UyiV9jEUdgAIn3Bm7BDzuCg/HnnBKD7nkB7qNlKnBzR6i5H23DHrK
pixTOUIOrnLwyQHYkwT3lT6mizP0BVrBM2u2VlbMLVdG1EOGrFpxGGu1eobQ/7xLvJ7g2+TBkpo7
MHVzAMWELmJoDcz/T433GMrzPKw1JP3b5qq+mDXHI083xzdaPSpisc9OqOhkqZ7xriMecJFnIeHY
0QGRezyQgTPRxXHi5Xl1E9rZsU6oFaQ2Cup4uH7LCYYGi73L92hTOVnqRtey3iD0CRWKmNbnLCxK
mfDy1lL3FyNry0Rrb2UFTuGh4HyjiuU2kObUMFpqVTiQC9CfoEkGx5h2zJeyn2mIxo5q7O9oGftM
1PwzCVgfD6S4W0aMkdTJS/QxO3PK8uHC1xG0gbqemn+HtqezT5yNB5RaTH1xrJnf7C72RDrA48Ix
NPWOZd0ASnMbhJ1Y5VvMC28/5p6mtxib4SZg1dOhINvkP9WUAQdAPrg1JjgwUqcQEffKXLO/GhlI
0tqOpSkLrxe6v5C4eIlFPe3XBnH5YFdaWUjC0RXw7EsDjAvFkagBlcA6mFMImDecXT9OCnVgMoj1
tP2XmNTrzHQ3Qa+4G0m99esxoc/w+DpfRoq25BVz9eVHKBz0k3vqvrDffCcCn/TXc3MZ7vGf6IjO
zRpioT7dywegvcTYzwfKNTSXlGtvGK7WWc4f5+NjYoah86xCkxueuo6ungAld9yt26psjd3Itr/P
MncH+dK9b7ehXdJhWkf1LBVhgicsxgIkfBt6vlZgmVNGGWV2pmU9em1n/mmr/3mmQx59NlkMTt9U
slfP2Mpg4+wtghvdZDFdj6phM1nAoUtapHtltcLZibRXM7HlF8ES6wDxQeG772cks20W3B373yns
1JF7t7X9mbMjBfZ2wMUb632uZzWGX4nspnbRFi33wiYceIgrTq9P5tqGrtktcOfz8MEZCzCSP8vl
x3P1gA5BEppasCv4mEzE4qjdT73YtOHt5uvXWRcnqccG+LFYCCwdaqj1TkC3GathYdw71tcvQUD+
sRZfOSXAz3bzaaAcTEEEy8T1CRvE7tAJp7Kj35hyWO7jnUFXIZFg2dMMZzxxi1GGpwqnxuNGzHr4
OtPOWS/i9ikYmimkwr8CbJCUP/qGnVeQyZqq1g7yRjOWuPTh47TspZb16+nuyBqpDMrPK9y7w50O
cYaqyPvVs7KBBhL9ipddG2digPyLoOTSW2ibqgoXGJ0v9nOLFJxWFnHEjeEqw6LkS9Vva2nQV/qO
Kb3bkyV1JOyj1tZaxPQ/cxXm/F2BjJwoO1agmVXU74sdwi0qr0V58jQWEXl8yW4beO2YsNVioK3A
mlQ05SsvbABcnL1oaAKmFyFwNAU1sovoFjNBRDjzstiCI91zAgfukr8KfTfIGTbrfm+R2PExGQ/L
a8L/wHepru9VG/cSpIPho3Qb5ClltzBi4Pdf4dwTjBCsTbSuccBtZ9GDgt9mRUDogRvHoJ9l+M5S
FbwdFAlwO+x1/IijDCFcN5MdfyH6cqxB4RIFq688cp1WN52Tk5cf7yP5rHez0pxh9V7v1Gt3nmV6
IvhzGF1Jib+ViVZe1jiPu6k0h18kfuHFj6qjk0FuV6UhC9uB1HbIw3sgmfSAJwGjoYliuSiztnS7
mP5a9uDluuwrvbT2lkzDjzOrzL7LoWSOF8ZTmX7gA/DNq7LTytj1VHpAo1at55PA88cy/ad20MjC
WAc4OT7zB4c/xaOR1pZ9J9pH5Luv4h1utVRvPA0tm/tyLJD4DHKZXVCQsowhjl8wDXI+8+2wZHTD
jWn6/ThIRKiI+jon1z/9Sh+sIeP/xXNvxbOqQhrvunHgWadoJy4ZnDMrzUhvBGbs36Cs/SfHfZ7B
87NEz8bzR/O0bm075PPQfwYFizBZ8GQobolLZ0EoiwwfUsC9E12Pt/DuMNtfNjyNNks86FU5CQAQ
X3mAFHKHzJDoWcRXr9Zt4a6WnHdBMWyjx59mdb76dUVcLG2sYW930nDulKEp+aHEyXU019917nGN
+S1vXbD/VObTDH/0NRT1ws22tOVlTZHXQBpK+VDZQQLbUj9QmEdwlyy5zkYR8n+jvaZTeC3QlNaX
4VtAoiYjGGS846n/DnPSoO8YaqotejUXSKHwID1GK1Zs8WqpBqBppaHYTgysGEc5zmvcw8DQr+6o
gqOu33n4p8E7Y5wnlKwHQLFndnkqu0/0NddCGckpg1N+3fXUDVbBVFTE3KacPQ25Wy68+ASY3e6s
BPg+YPguHS6b9La4QNCzbDTB10Gm0SSn7b29PCmjNmqYQl9Lwo/xar9mXozXbKddwNXe06w7/wXp
IOetl17SoQb7AVS7LNbrDsuVKNzBXycnLwD6u6sF7uT5ugshwVn8sJEBWOlxxB/4MtF39A9ZD/SC
njPOyLU9gau17U7J5nlF2ST4Fed0DNf+mUtcpyPxX12jNmVt0tT0DiYeLrKEp/Ex4cyaD+Jss/47
chxTjWI48o9BHQXZSH6RA14ZhMOG1iUZrroJmHA0efmF+WzAkgz71ZV6xFH6Lh1BHs5BEIa7nSFo
LotZNubk3+Q6uFvHDmkHE+GzF4pqxPbL10I3/wqP5XyggTEq2Eev15GUpXLpFQBLsgndipMsc6Q5
GYDlswATkUyl5g0MQxQSyqGO/TXQs7fBYaU7Hv6jiK06G7XIwRlOZsUkH6cPGKM1GniwbCAtlTx5
XZ5QU7bYlV+jn68OMeNA/BVxKYCxDQSM7+KWsVJq2sWQc/Hum0BUVqSdrmPZwYW+LmaznanTl9ON
W9ltxmu/RadJbNpcuY/WWNQBtnr7BeG0VQhaaW5FhZG6EmbRwoDoj1xgxI9Ts1GXe2vBrXjXjjiy
WFBTkJc+WloponNbGyj5w9RxpIWnB7EJK94zIgmcar/tuuMA3hRoO+c+EuL/033JNrEk06z/6cfD
3V7mvrJa+YvIRDBjq7qQE2pXpMTCcp4w8QxTIScIga2dIceM0bLa1o4EqDcuPCYMlsl7bNpMxwgC
WpotYqyiZ5fmdxkfUyFiKl7PqnceBZzLDZtRLFwEppRjvGVly1Zjdrt/sfeUxMzegnV862kOAIIx
Q8Fxoz+M+cQ2CcthAKdQABIjvErWS9t59KFb9aZ8Wql5On5nnOGTX82f0givW8vRGo90Umy6LTGJ
9iQf1J85rkXIwtMgd3wBEqw7QpATNaxznUO2VR0p+0ZYDxUtPwHTnt9U2x3NNMymdYnHNglU87lA
8t+xlBU9U+IUEPSlyLi3IXX5GjHlahGNHXIQfr4vJi3SSSa1jM8vKO6HLuxhDnX2uM3MmeG6bx/1
xjWpsWQyL5meG+RAcKtpVSOAccK2109UPhfB8ghG264PIKfq/ZcTIj5OdDHcsNm5HJ73KBtlbaS5
XoY278FZuTdbML53aM4wwRTucEBkILos+pbIrPhPCK5kkkh0xzcOmVfOeB3f1uICVh/mUvcrxgqD
a+mFy6R+b3Lx5bX5YsFhx0qoObdgGnrapUUunmM7F4Y6/9yNp3/EXhSc4RQF0x4daatkK/goE8UG
TqKh33K58dP2CLZ9D14s4wZe0MDU+t/0CVTllMG5P9cO4NjSFup8xSJj8iIw/byB5xJbpIQrC6MK
qO8i92YOQSqgK0en5ukhHtTaNEE2/S1E/nIijoncotJDhnTuzJ5Cd1KN7JgDYz1kQbcOpJXk+pL2
J+rHqN4kVbPwScKLOE3DIvTY7zH8IWxu/vMHTE37wNIRdPMXyWzJmQZTafd52B3BEzmh5OaSbVsU
ocQspztOFxD5f+ViJj+IvZQ5ORC3NHuAZBM7nFxbKj5V1pTHK9oQQbhT8PvzYXe23D0KQVc1WhVl
BSmQVdsOlymdochr/UxnokfyvgdJgaRGO1sj+zdN/76XZGc+U+ZLuvHBxBCIf7ZJakPQMPO3DU0Q
Nr9d4mAwLqr3TR7w18giWQAjy9nB7TyllDr/wmlUld0wDIZZEIl7os59Da0rWLrhXV/c84GdVvby
+a3HHojyRGrnHThVLR5fHL98gtdLl0M5WFpNe9MNF8AxwiikVVyt2Jgrtt+asVK7J61RQU/qzaL8
gGpcZnIJCXRNuxr7Bm724Jv7e5oD86nLWPvHxSyoY1GBIFUl7bo1fqG8n3QSvAjbCIxxli3rK2Wo
kyPNnsbL7cvpNeaRcs4OjUXZ32X6zsF/eqrDMABpLUaHBhaTh0rEJ1QqJnhTR+ERv7TID2wqXcG/
HKtM2AIO/rsLRvPxmuQ/56DPAKBYTc/PIpOL1tNchfXcAR84QV9qOi0iLRT9jMDO11OTrbBFQMuj
5GbGrWh00Aww4+mRNAw1HafoJI/s+Q3h/KlBOP2TnAUMjM0cQOYokxO3mt48hq40Z+5PrHY6Vb+3
g9RiEZoicdDTBuYh/ERz4bWx1pz2y6mJweXHDg2yqeFGcYqmClFcnlr9et2YxK75O0FOioMyiHTs
QCmpO8PaaIS4hR7gqdFXoL7TT6ygfVbpaKJg7WGFtpMxElF8zOCE7S61LZMoIbmSie9446NbpO6h
cg8rMLq2Qlj9qEWgmAb1WTu84OOTPhXYTf0vbC9KK/kJN6RshyW/xh0YEsqTxH9qMMhBXiz8iAHC
Ho2A3Owi4aCwD9WrNs82MXXpge6bPkGov2i/BEIIUW3nnXmfQV9m9cAMpfYyRxqJrJtyVXTf6DhA
eTbIqgtx6E9iSEC8HCFufjASQKneP/47kGPTmS8sp2xlIYCYCIjK+sctXXxbgVzZ4DUkuE/otcGj
+SYaFJLTKpoRoEHprtjyknYZFyeIrX+YWAacPh1chC8flsJrQbOB3SlHSwJ1E7GdtTTOlMSAq/Uy
67ID3Y/buua4ywwlVRJ/xIBmElr97QJ+vCfPwISW1jFioc/WJa4PDVx3MbXlfsJ3Xi37MptrLtMU
ss8myMU3mrdNjpJjufDkDUifT9fi6a035vFdxJffHWctkPmIJvD8Qgsz2VzAtvIuDtMe2FdMjXGe
fNWbzAKYbz+1lZA6AqhX4yQ+nYS+y32VAdxhpq4JIk1x5snXhuGfnU2sGJddz4j9MPXaBer4MpQr
4fFKSdBsJ8NfaCDxpeaDZF9L3ZrFLLus9JEUPPWKzSgvNU2lDYXw5G4q/HzwvqZEqsBlz3Z1bjUf
cUOQ/lvc6GXygF4M0+57T7UYjKUl9QPvxa6uchOEfVqFgX6TX/BWiW8qfLVXJLV7NoF4Zjv8ibp5
jZWuNbclTj1BJdLU6b8/R08gcHjQtJ5zxVLHFuLgZfM031XEebI/QTLVd5FPD8eSqEDzxpC+Vujg
P0DY/oAkJUJiWxJCeJJ1BCrn7OCmM7c7+d1/TowXtW9bm0/huTOvjnkG9krNgKBg6MJTdpnus8ll
nYakN6v3PTaVp8olHFeYxLV9E/h0n1fNbsm1YsE1ay5RxmzQ28CHBH7WaqTgd/dNwhKqp/raOQpT
eEiIrnTXJbDvtueD1jA2jf19EFcNAiRkw19A8A0BkVLcl9HA5/VnsRwPabXXAZBmqNKxc90NyDWF
nEQZHVDNIMXxW1XMGOtNnl6ceSInYPplRGcjYM0Uyhkcs43lcfG1EksgMbv1Pfr4pQa56iFqWVFP
l5J+eCNVOnkryxDnSb2MISvaqmwAwH9rsAM5nOYESJu96GBNWsYDFCprNhlYGTBJPCA8HJvYTfwF
UE9HmNaM4MUjQCuUKxM+DxbDEv9yI81YRQUJIL8CFdM62C2Q6OH6DPuUDY6bf4fauyeFB7168eap
+M4AMl/1veIufv+S8fh8KAl+D4cuf5VOH7c1NGXXi0trO2TO3+fcTDk8onomNmYs9bsbBm/Utkyq
b+TCOotOFu4jy8da/gIEPo0oVVLgmgUtchq6ADxDSpO9uvTTZCTTnNw9VxiImTH5wEu9mMFhL2Ss
TLUrUPUC1bE6UMz2EsjppfXjPb8kDKMoKuxJILVaEaImO1/w2AWVxBgJsqFP844zt8aqPwdj6TMV
IJ8ZE6GAPH8+KDIYRljcYs3NOXhkOSAntwUZzkvQ2FDJh1mIJYCxo5nTB8NnFCojlSL/6v8IhNQ8
IevIjOshPHXV9p+yPK/vO9EpVb6yNkjkHPDjAzYqqzcKXVSWsh6lvXtthy4Wont5jVAaIfb+zt2Z
2b9YdxEES7O94L/sWnGBNQWq52NFTdF8RusPTsgSKezriUBBNUFsbLxLDunhJF/TbCPG+NX69cdm
ci76sA3hcUvyaQzl17qvLlGrqbi3n7bVjegcGPxiGQIfjvg5I8TPBM3bYw441Ge04LB3ZtxAA71K
ZDehzxsBsnVFlitDipJ6CHW9B9NEhWy+3tv7aiFK45KnOudHrt2r5No9LXn8yO8GAcJRX4xG40sc
J97Is3gCFEAoXU6z8+jVFA4xXrem7CS3hnY4beySOppk87/WMzJe+t+L7z/TWo6of/ztLqT+Tr8M
X3aoRJsIYocs3DcW9DS2v/HzovdpQcMl7kbKzyelSw5QxNcE/vXmKSIzWN4H3Xhrkuraqs/sS5dv
yySkwktuYbLGGv47PpCrbIcwk1ssoHufJyHL2VI4S7vmARn1he744bcvsbGvCTjzCZlSEiU3rZqM
aRkyETQ5kxaszkBytVKjg+tJKbjRuUBV2arOCKmpgpXeozvMoj5kEJp4rPgd1UBS7l+AXJ98KlkS
yWzGgTYiXFD+hB0eeRS+x/krvvXNcAzaahCsYPfAmLUVK3Rhp3pcOwrQn/yYga1HSpunGfMRjwQx
AX14slAHPqE9ijDwgN0qFQ4phT5KMWUa9p56X50B8sQLc2WnzwPFuu+b6e3kHaomrnSa9huXuS76
sCzVhsq+y3oIkBukr8tO6jgJR8XTzlMbdG+ygjFQYPaDQh2aNt9UJpLrgbyRxCt/BeOIL7PT0Eha
Rg6jYWVkI2dH1ZomZx0dQmU0ZkHEtIMGjgNa/gPaTHxhyrwy06KkbhcYR5Uqn6rlZOShO7WGs/l5
stps4B9TT3WTNPiL5eH+ssB6dp5ZmN2LxCNLzsew7Rca0IgAQp6/X08+vTTfpzq0hkaPfCzMDzgX
rLGNPXJqeUXqL4X1bGRV9Uv2kgyhqv9KEplVJ3C3k0pUdvLlh2gygynl2Aracg7WGEIvXqTUNGtw
LesdLbO9k9EQ6dQiiEhzCM+uCaVJyiVHu9aYprp3DW0L+vw+obz5sQ5cuHOqqgeemFzV9anpv0hz
GVY9dza/0OZHNCTWh0um8/cgj9VPhsM+CcpD49qV1dh6oRM2TdEPV2tp/DLUwLgngC2rn6bndZbT
Lykr/lBW6UkC37lcVT3RAbSjj0byfkzXySdvX4DnUT5dJuFegcGMtUz11/96nsHhUuyWHoOozHGd
vFqqpAXQ/q00yRvoZ/q4IJ9AZNgklrwAd3FU+OPwkajFq6ToAAJUyLaCoe9c/V4R8MO1RPoepQvc
RM/AZnpmIW71oFUz/t4IQ6NbRbb/myUFgcw5VV30a0wDdE8w5SsBys9yANuRx8hlHmQM+IOgFCyP
iBBePSlVBJ1quB0D/WUFt2vup7LE25WHvcYlMHSIEQzDcDig9Up6SbL7qChnynIN4i7YDcX63cFQ
+2L+j2fk9bSvj/ozzTdu8NHFf0eNTR8w9nuNtzGeZYknunCjXvIdLTMD6+SMpVnIUb2unQX/HQcS
hca/MtpHP0LzqbvWXTn4vy9naHcIw3KdTdXIyiYOBeRtxu5pVI5w9/QHrWk0AthfcCdSEHdz+dae
NcQ17O96Qe05aG8KP0u5oW0CQORts8hmcDbu1w4+TLl3Kd2oDODSvdYe1TJbUvryy8hH91KZnQPB
JAQh++9P8NIWruqmiOfsrorbbY3S4Y+76JxabOg7UKMqcxppOVaUYHyZSDBuCdDQiiD61QjJGGvI
w3CrdaTN2JdygYgi75YUgau0Fwbsqd/SyAEaDXps+F2A6nyuhB5iaQbgs5/pji4ilxiZXBcAL2c1
/f/mWx6rGsprRoqqEdJVbE6JAsrDvpjOOboboDctvEituO2JfNWTiiJ+InXm9mIPUQaXBredXeWD
qeNE4cs5zchOR+ARR3ABjdA0W6cM2BUSbrtjEltyjwmpqZDlhP6qSfLNKBZC7WakG9J1SLCPFNig
X6gLcUjfTMTV/GbTzzYh1tlJ5t3gTgPqMe/ww4Tqd+6O5ABg94GXOSYPEtDuk9QS3oOjoKYCGACw
CbPDLmuUthtIvLSiMyJ9ee8tBEpzQ62fRnggzBGyf8zC3GVj68ZDE07GLTrRtK0YPLBIr9zrtP93
xCLY4ddcMHqfrhhNWOotwCeQE/2RRrZpJwaJ72xBCQD5TwTqOftYdPobHYDjrFY6x5uC4Him7OSF
EClQ0veZ52f2uBZI0FCqJaiJ2qjCBtQi2X2bEpQFk+sFejLUl70KasB4fJ4htF+teNZ3Qb+YW7SL
Z0fYjbCZ9JRghsd7pkV8xWhL7yrK0KYI1TKqQqYWqP6cD1bB2Y+1Fk1uhA08IBD/t25CX5rZiZUI
y52a2bBqO3YGT5v5fRsYLYdvriFIagzJbU7xRswjekFQBFhIGLq7DMp0xdW5GAskCGp//MOKSLzM
x7Z+oF+WlWBb9Wt6S7u5nUv/30PGyfr8o3BuzaiGTTTmzdxTd+LBTwiVjGzd2S8aLMVIOZ2cMKJm
DaNV57YDRgQDe5e9VVMOoR6v1Gnq9wK8le2S787cKVLgNF+9G5ul2RQoI7EUEVod3KLcKS/h6e8O
QXNhcStdgGjWky3QgnrIboDlAnrVUJ3UHDJ42mB5Lh2y2yJ1kEeAdKCmlcT8XdJypusq1JvM7ay3
bGYjrMhdiqq/5Ndx4N0hlYrelfAXims1Awg42kb80e0fiY6Pmj4zVSL+DbNU1nQljfMUx2iboBec
ymkmjWQvzoyW4FDoDSr2y2XjosCFJq/TRFD8pgWikpjhcvOiYEcWsqfjl0MDuzVp+hwnqlE4luYR
83HrqJLVtsk9WhtE/ItVMKIE/prV2pIiDHxxlmMOuBUY/BIkkQYt8pfM2vgLKmcDZKui42wzXvll
AnMELVBW3KyEDuN5jL2JCLVtkGaBq2/qoUcMTC1stuHIk9PBwkRqSBNf9FuL+/ZxZuE0JyRDvQkD
tKonDD3CHJWr8QhkchTolH78aPWEu6fm2937Y3oDo8PDzAyfjKtZn2pUS/3eGhc92E2LQB4WM2qA
Bn2C+oynIBD3RcFL6g13Swu5cV5XmTiB7WhNRpHdWHcRvmKlb3CPe2cn8+jRhBxlxGL/ckbSkQD7
W4rKXyk4o79o9dPLJl5NNky78i0WkG9dza3Y1Z5yc6uf470hpJB16nsx9znktWfTviByz6hVdQaM
IeCd/QrgfqFk6Xlul2k1D/YQMcIWT98nNSwQx3A2Ot88PljgyePvXLQrvw+caC5OhujJJJvplcZT
TWi+LvYszPoOluCWDx/rXNgnPT+HSjYdSFtUiSil0Ut991AE8EN70IUjOS3x4xSQmw5x3UO/PwEm
R0cadzMga3Uo2rQynQ07yhNyCed567Y15tqf8N/aFV/9WrDyMbHl7DGBK3LlRM7T1Qm3YPcX29Fw
mgQ1gwwAWNCMZ8P2+ycoRcmQxrpU4sXgNaXtSzj7Y2xC/BQAsNnNsDg/3AMzdTn6ZhAtD5QlsWLt
aeIZ5JxSa3uriI6dXlBi/Gkdo5ULb+1WOBkN5hR+Fvp9ASiRZmYcXRbZXd0/cAg85RAUWXq3iSuw
ioLtwEXc/lfEQ5qqlozjLobSqCL+7rg8m6Z8mWANwkAw+N9Cnzv2Y5BYfN8AoL273ScFgl3rZN7M
kwtdG122Mq9pHyjdTq6sXOilW88P4zaL7WeG+dQILRTieKlsY7LeiCipbhGkcY0oF2mZH+eRWbvN
eok5XGoKh8F7N8sNm9tU4GluwCCGZ+zr0aDJAuoykzUXoajJKQ5MHZ/J3HrPUTH+zAG+oiSObUFH
iAyCT4GAygnsEeNeRMkngOfgzb1vfCfBxLpRNdQ+Lkr+xW0qexbzPCf9xVR9MhjcpEqc+M+UDedu
gxDjTvA4EGK06NpxiAYRgl3rtp6ntGSPd0gMzl0z95mZ7hs3KGMxLgZCuF2sjTjcB8xczRN1KIxT
lm+WMVzhvHWgtuECAg9viGUVcNQbe+hFA6D9dEeMkfma+4/Gm/JD14/sI/SL/QYx4lS/C+RhsBLv
PVUqmtxwh5tG1/7brujZSmKAZMwZL4NN/V3Yi7yONjG0hjPp0xZ7p+UMkRg4qTr5YX8/mqp0bLI/
1fX+ma07GfWopPNO8HNtSmvaNh1AobzaqLOtrEHqbTNoBr83xD+LIEGy0YVjYJXyPmTeyVgvPjDX
4MUhrb/e8tN1FiQzwYgUH6r1yBj3/Bv6DHuco47GZYKTDn8V7swPcG5kGKpj3X1nrMWPsHebR8kM
Im2WZgv27o8il4YWRD9ocImUc5IUERbMBrUoMN+Kg7uc+Dzbmw2Y6noQikxVYMeODuIhIh71lheI
NyndAPPt9bBm3f0YFh08Kh6rmL4zpaJxWv/dpU5V35L0gLkaGnX64dOpK+x+7a3QKf2eNa2qRWad
PCuK1gbwRpTroYPeNcRNc9mnaDyQI9TtJfnJMKVeLdLRItlAPFl+9I04a3lYhaTPCWCcPhw2+rGW
/IfZjZahBrtdxovEAulHg0MnrozI9a+ZiWwmGVHXFrNSlqm6HZ7hilR/+zZaHJ8BHxiDVyw+3CJx
e7zrER545jJ5ul+cgq9Gf6DP0hhBxyz5IMttAtxTC8s4+4WoF5KQUcoGbw7lua9Wpk13Tkk9YvEC
MsVfZq7dfUNpHfE8bXGsLmz3wZsdGIBuOMSU5i1SqgZ52JvKWO2nfzmE4HpcZV6/8TVDQu0RJFXp
XSdm7NewmIwcDojP8E0clxDFhINkbSELnY04VLD7ZfSxSmNgRCJuToY+I492K/eEVOeaKcgi3H3a
rKvXAPbuDfoS5YJmdIfl4KWHbkhaAEgDAklct4ZxcuPFTOjWY7WbV5gLyXJJ9wIBcwFfKas80lHx
8J6Cv4KxsHY32AoayldQdwq6xEjv4Q4m0jIYNvHDn8w86V5H7SiTzyMLsprsSVW6K722KVO8Jx1k
aRKahY6shBOGHyb4eCMG7cHuC/lEW5yDSl1OCeWCKfd5cvjQDyFZVlJPn+H6DRmS+DE5bLDW0b79
ks4v4A0op9P60GjQJXt1hO+1m4OrgQUnfkdvYi2MBN2QtmqFHco7dq8yQrzEdYc7Ea36glSFcMqR
Ij5WY6hPWGkvzR6tC/+PewSOazWOHNLFp0YPLUqbhKThb62HGWXSoQKuD4LShoj7AeEOMWxoR2Pj
lMO8yZoPF2VS4oB1itvrOdJTrZ4Yy0EexAZilHGgsKDF1NW06Qf5cNwRRZ/tAeMsOdgLIYu4mdGD
yxsH1W8rl+kL7rAb2v70oSCt9MzoavE36iTJND3MNGnKTehGPwUl89hEp3WisAGUfubskQ51QWHT
OaZ2BxwtbQhy4Qmi3+B6zpJKWnHdhXSesEjLrOGvv1DEAc+8hx+xQzVsDW1+41/afhgilZ4MNbXz
1sINCFTq5UGIhL4dJJADJes9E6G+4xuKsLppxsHFEkLoUr0nEpcGa2xrupcd7I/Qi+jkPGqpf9Ib
Re+wn2Hsd8QLN/bk5g7x2AeayAGM6HFXDSjSY+CXzEZYI/XMAvKKszgkEdR6DEqU4Ef7bUN0D5WE
CnzZ35PaD4pkFcSFbAMxO+oRBEDJ0K31aDSDNVEj2BYqkCeldDdzhkDGrJwJa64NSvU1ZkrkvJvi
pkQ2CsLqF/B1WfL3ZDiNconmCkx0qFHb8QgrpmOv9O38z3b+LCgci6YNxbdgLG5hLL6lIp4pe9G7
9Uo9ag9UyuasTi2zSmJyDg5EwoeBB3a+vUFnj0fSI0B6PugwLcrNSu5CXurODRaGb90bE9BoA3HN
LYm1STD9l679sMqPLdcrIKeOTbAc7uv5IfH6eJkUZu9zDOJR27bsUkpC65m80w87XhGMDirmyjs0
KuoPGppMn1975udSFIa0n/6QpIslAFbBtYwuLbl/xCc4JzEMROQcIeMWUq6ki09elyI/MqcPgXOZ
2c+P1y0F6gfFHO54Dy7b2cIdh4pv1LD/KM5JYM0nfBnl/Ng6XPqUhHv02eYYDMojB0mPzUkJu/Gj
Pjsg5ehE97vjwffP2PjTY0ReeaMQvG2MVQNRvNMr4cFhqkWZTbablPlZtDpQ/RhfNu8ap3PVvvrh
HnSZC2ucJRwIAv9acvbwNRMfSfDUVqd49jY1heToNrEB9jiZPXOEK9rFN6B4MEI7Z/i23qck3R68
MwzjxfBXplJ+PlxEhOqg6Aq3Ey62XXaeH9dedpXb/smd5k4otgLu1Fa0SA5Dj6poZGwNbZjS65gs
krLelBVh9X14dn7ktFlBXhZctGiHXjgUhaj9XcVay4uA+2bv6R/m/sen3xMbWbeNHJF9/GxSnJ4X
iOeSJG6xQzwSHDV6LknmrgEytIM69yvB2GO5+klTlXDJ7r5bw96Lz9yZDUBDsLku3imqEW0ByqHC
lkEkLLb+fPIi046vgNQW78s6uyQVm2sXqotEkDFEjifRc1xhCX3Sq2wR2AVvD/uFr7ri/K2duat8
Xc5uqqi8H6g7i938RuqDSEbNP3OOFGDC4qvYi2aL28laRvRw/Mp7dSS4QM525RREclh38KbJ/ntR
7JRuk1q5N5LKxHIctqOE0Kn8aCuX74XtS7suv+5zayDSHXoM5gQNDFtaaRgLk39onCS1MwvE9dV7
73ttdXCCPqaQwuPiLcM9HVaCYkE5rgBv1/4z+kCM7cbFVLfsFrNdXJnvF3LShQyp+qEC35NXf1nr
Vykf4MFrICGcYZxijnLJ2jB/YuxDogzH3x4KfRebN0SpQuFuZ7mAYzlIQU+4MyTofjAunoexwv9T
PuZzEegK94U7JjZzcaIq6j0SV/ATH8mG7OyNaarLAc8lnG7UFt67ijnCrKJJabL/bgD4w9+ggved
E+O3WICuL3bvxFTbYk0wVxTbURW8zBKCmioaTMZ2ImzBydvEwmZYTmej9tqIQgKxXvmQ/fx399ZE
eqqL/PFg2h+w6vX0NNZXS0m9ae/lqVpj28h8UINkYWKALWh7MCV2WNiC9qy+ZDtj72FqQRjLP+VX
kd/NwqFd93BFpDxqABFGGaG2vr9itGpq4SNt/RbtPiLM07ATdW0lANZgPL39+oC0RmPr/euSQ21g
yAWMtr5LIVxId44cR9ruZ41eTYfG3NbK8Z/V36gWBsEPzIQ5DLl4r+yuUfrUApUF1Q1KIzkwHCIF
NmFj9oiYVRPCrYKqbY8AWCsgldo5pEempzsde22KN8PEnNwtGG4wN1eTVM3Ka/x8fieLvT5j+S+I
SpdqO3BqS8WP6Lh3enSeNNL+xzJnk4OjMw9oRzS6Nxymvfq0oOVwm36yy6ZM1nkc/dUzOdMo/PDs
8dkAOW8Nnw3ye9FflMOXChdueRC9hgY0bduFdI5wZtWgYvcMN/M4xgq7+VKep5nStTPJVBPk6U9e
h7T68YYjXfGzfhCpsQmADacDbBs7x8n9KDvc5AhkDY9ihej94rBGfIOD2t3OL+bC4TB2Tv3WxVZe
so8uDZ9AEfjgRcEiJqLd154jI9ve5WE9fkucQqpYCMkJ0UVq3MiqpkFSMv8pmL4asqHGTS3O7li0
JDk6PAiqVUZ96S5E8DYbL/csoo81Q2AYobbFT76obM+d1lzrcONMZfdafJMJgS9TsAUPUwjPh+s0
ba1gTARLjGGoCdbT+NjcO3Xe6qHgIRJLUAOU4GwmBRaPgT+mViSbbGJopO75hI/MEdGajOcUgLlP
mu61FYQLJzHEmB3OINVWVIfKRQCnw1lY+oGMpaDu+5EoQ3+lA12ZrBXd2KE9tcPPKwEJB6uC7RbC
/tHiS+zXcVml1bvTL2nuYVzMLWfhvQGzRxZxs6FOWEx06HiMRcauIB4WmJ83t5+H60vXEtQyDp5q
5Ff4YtoTtJ0hkd6dmvtBD1RJ0GH5MUxXVUcWAL4WX/w23ox84hO9Dx/QX/Q3JhmavOCMRxv7J8ul
NCSWqGPk40to/cQiJEVxlmWctZlRCI0BXT0yT2lr/lOV6w1DH/4D1rEK4JjuDcvIyFO5GC10ETnc
8I9IlN2triZKuLm5b+ZAU2F/Mp4qvqQh/cWxf36ZF9U2aNLsyiz0712zi1m+B3pT6pVz8N2ztfLS
HWQ1BpfN7EQ2+eRUTE8O3N8CQbDP5oYqD+U6Xo3Q7+nY7XwcjtccSiF2K4fwH00Ri73tGoMe0DHr
A/IVjgW+miqSFt8aGJEBQ/rgak/xqU6c52/xc5LiRgvp3oXb2S3AKreRGEz8m911BovcfwjIBTp0
8ATd2tPmO/N2NCJ/gL9+U8QDpjnBQX0wIfR6x4s6rIYM/gSX9+tDnw9Qb3p4FH0zt5beevOQ/1NN
gzClbnAioo/8lfA7KsNBs7KAdEy0bqrOg7Vy29xsi0cWSNBz4DJ+lBangC61O+ilqiZJzJxeSr1l
Yuzt5HksNmctKOCyhYnejtB0R9AM4yAY2NPqTT3Vz6PofIU8AxC5PgBAFHa97Lrp3uE41AFoOEu8
PG95IikBeBxGnZbfhLoaLY3y5ktzUVzKw0buRFLrMx/HwYWF/HnG0LVGYoyhyfRgZg/L+o7npVGt
sdZE3Ag4TAsKEfc5BFpqNNsXMVX8JZt4Y4ozClfkj7N2njaFdzEn0++/AueR1xHRnRxsS8nwZXiy
Pm6EtHQPcMzmg4daDLvp0mWVO+OezN7+oblln9NP3XvGer4iR7/o2d9TGJc13684Gg829FnI5fyI
rXs7sNk6+xZktZpGI1/Fs/9yGSOFUGo1qJ/L4YAxW1+g1Z/C/9OBfaYWialLhBHFnb+KlMHhMT+D
MOKYR1Hg3B4brwEfPcMOVZJhlzEfjFvNfbO6W4HS2fqvXEd2w88clWYcaijamg25YeiD/rcawHPA
+xNdVMcg4jBvW4gGt6nmE+tOcBgCwuh6LN4Kqnhk2gwwlaTYQHqGpm0L/jgTN3mbjMolCLOIJdn0
kpl9QPo6ancnBao1+Q9eRV6X/aLwF83Aduw53fJSi4lyr++PqM2M7QhJE5uA8kQo9aYgTcQSZPce
VZPoyy0jgFYhDnWUBXkL/k/xfKX7qhe2a9hfTVo1HQkERgGRe4xsZrUO2P2lXa1BHrZ9M7+9HOyf
nzEiLvVHCvfWNEs27k30pSsZNCUwgZJTgLa6hOCm5BjdvIGQ2sktBODYyCWahL6CV6/ctPLgcsrW
/iQekfkbN8LRCqAdYlz/sQC8bPpcXwKB+6Xcg/nUa4LH+SNLibQD9LoB9AKP2KFYIIdP0vDZUGdp
b6mXGbuznGDQCHMh4M+MX1bwxxC09ZqLTizRL5ECE3WKfnr2G5aYRM6tKFGDIzj2P3H7ocM53Tzo
2s4Cbke/Elvu6dU6udcjJDvVFnsA7UXLAIi6TgLG2LGCPndH+ttTeB21iTaL+wawv2owwcz+QJE6
CIazM8UmIewK/fZFpy6EFq2092wHifz2mmreNP5wWQG03GG0bKQdChbPpFLWKRSewXYbaH5yrHFh
4u43FNQEQFUR8AB9Cvac2Bt2i51gsQX3fhsfBZvRnBzbXPs6CWLIHn9cMx9A4ohid8ephGmmDM5h
2Z6KKxMlHW9hm/DXILHHd7E/bCmAdD6FeNcitX2uGEOn210SpvKXwuVQYOgQnKeK7w0M089VNrRp
MhyHFdNEev7e9PTrr7GrjnsvuqhT9R59mzhUIR6K0Gjr+kb9otXVrNwAoUTGGbPL7xQr4qDo9U5r
0ZNkI8SK4d59GDNeKlJD4eYnYD0zJ23YDMzHL1qoagsrZ0LzWu4IXBycoHj6GKeGdrhx5Xo9u5KZ
qkc8wKB7VuiWTe3sPLgKGLnXj78fx+SqCmrYAGla4IfxjHiAXCUfBouw7yJ64PlYaWO3TdV0Mz33
Qp+AMlSxZlcpzxSImeaU81+0TNbkw0LMtdErOo9DUCeD/VO3B6OTqDaYRfEKCeUZ2jiX2jq+BojF
MbEl3cH3k/pLqcSO4J5zWolaoPGJEiX3JhjUFA1P1aLLow3KRK+IfcILIuoY5aAm9Ua6fjDWDMnk
VTXedurNFetVkM4lXhTIk+XhqierZQ+UvvyUQ2NCvOQOivdpoFvorp1k6mgJiPT432Pw6sZr5Vg3
IR798H8xY1wLGAbQBy/xlSICLPV1W+Swbzrq9Wuw7C4Fnq2IljRyXX+uLoRuPJpCIxP4HzN9wEtl
NK+tjpC1WkS+9dsjo68GIjQfh25pMgfs/0SKs/YkWLOabnj56hcA3LwA2yJuYhkRl5yxNKCTEvM+
ywueROM9Pqt1LnGtYla9eCXMVpC3Jzc7UtVlIHP0ITdjGr0oqygAJXH9x9ZsYZy+Faxjfmzypc10
ukO8Yj3qJAnd40MUyOcAzvMSpGh7fuVh0xhOT7qpp9sstNtOUULGGatHuv51CP7bmpWG4ovqMj2f
BQFXS2dSNSBQEFr+ZouGH5jLDf76YWjtDBqPRIgn4EaO6vyld7jW2t7tQwoDfDRVNy87n/ParZ7L
Vtd+gzqHeteB3eOsI+5DCf1JzZLZSsxMdNv1dDD9eKx7tGRVY5tp82fwiWr+8IjhulrcMY/k4256
RmMZnrZhz0OjBPxM8Qiy9pzIwNpsPMqVZqWhUBoekpMOiWAQ45lH7xwuLirmF6ku9b4ZOHXdI78m
81VZCNkU0Qy/eJiuz56U6AklrPr3wdQzXgUWYhtBXTNEV1RFmnqZaOUzv2HbdacltsPbsDWlEK9F
YaJD0r7TkRcUxITunEiM2E3rf9Jr+HUrlhZM+Hr3Nnop8KsXqc2s6pFVb0wMTvrtyRe6HabKIh3p
9h/s937qqhG1cYT+thJnQQgihEvKGpmcR1WbkWhUxMUhZhwzjO2RgBDl1hAQA3AZbNmrkZYFOnyg
6DCBZCUe+VFMZbaTcrcOuCOEjr0be4dXznQEiS9kAyum6tABIRpo6wtdIrDbsHaWMYKf0LD1TuDG
Q5J/wucZwpfexgDlKs7bA5Cbq9s2pGpvkg13oGMJmq7H9zd8ZuA9VyNmp7px1+xwYt+bhOnxXoyP
3VWk+PSyScdmmdDPgTCklWSN2EbVcVtvh8vPJ2qYbIj2G3we+v+08JdXPnawwqv5bATvHu9DWN0k
g3R6MFIWXO7nY3BEs55Rbh9KlEqFdl/YizNCpIQZ1PAfKy5VNNZSYAofgspk6ILFDjT3zrJ0B3AK
7uSMWeLrRXBBm7wHUFMxIfMkWGAbUXGq9RdcF/c24aILYHqz17NstEol5yQtg57WSPzyA6ueVEhC
jA10o4I2OMu/36GFxwMQ8rBsQcvN6KZfHvNvxUXO0aJx/eoTBX3GA5SrUissHZuEnoN1Cw5nIcRR
RnuIQ9RZpbM0io+UQA5VSWWHyKA/crRKmz/L+4rHYacGMQ6LtdFpf/z+TafGWAdF+fS38Mf6br8u
sPfZ2vAJdqEwmzSwB7ii8JF9A35LYI18EKaTCvgHmqpuMwq7hy+O3oJGHPGDLOQ9fRAE/R4O2fWM
OW0CuJrBY8jUULYsr55lS5/8UiY80xjxleRAo9FHQ4ejefeMn3ye8fBd2IPZxN3sFwz9M0N4eM0J
w4ghH1R/C7zQzyJXDOqKPOWo97MIgp+Uzs8VZp4V+AT1x+OjiuDw7ISzicTZmRZ/1e7i06DrrNDG
+Mr96PMQyzqC/jAX5t++qE9I/VnmUXVoWyIZHpMddoSnd1Uw/wuuRXgJpw2lJQVCzzCa/GNdzPqE
C55owFNchwqlq7B9FOWxzRFQWwPABECD8bXzo2NbOvDCcoA7nhZT9iFW4cO7kVgWBLrmgDuvIEZ8
ajWmfpKfSX7D5Lt20XZSFV84uf7b+KV587ROMzP4fbuLmh9PVf1W+Fba3C2DLVgRGBIxFU1HUEFv
QyBIWKQM5Qi/8j5rQ8kvw9aYZKidpMRi9Z9HJXvt6nHnpwRX0YRYlMvPZlv00fA56ML/uShojRlk
IOoKpFlz5qnREWjAv+C0t3RznxMqXf5kSjedFyI6fnfgQtNU0b2U/J1M5Wc/cOP/El6aQCZ2ohPa
ZfCvTyNaV6bUuPjCsk/iNpphuSrX9NOUFZrd2Wi+gK6ypGqH9zR3VLxwLOwj1oTBWZOLxy1AmL1/
HOA1GYjGCAb+hNcGyNqQAsh2kV82uccq2d4sg/DxoDFQcavl30XNBwwueGWPaQnNNDDf7+1OxFJH
KBlav8fNmh+5SyZFvV+pBBfe6st1kJiH5drQXsLTWvZ8w4AozB5Gwtdtr8i9tk4yyrXPA4mO3RM0
m2JLNdFqLprUX1q4gQprDQTx3X9cy9vJwwHwQzZt5llpUBUIZOL1xNbvf/fpqtXl5gWloCKWyYs/
8EG8lct8TMeYerWhXMPGZ/6OLgHXxV4eyaRJOhDx/fopkWzgqRdInJBwWdH7zfhYRdLf/2uAGODx
nxGZdwYS8+Eni9PPX8cdc0dMv+xQMvpL8143KWRCr9bIhodPYhCg1aDtPJWpxFEv5/XperJb5Hzj
IETBs8doyhYU0uzm4IpEwvAcLJHz8WJEjbEH+cDptqU9FG6SKRa10FfI41YesnQNADoqGu2vYQmk
n0KVT5wJiiEvrr6iZKSEKucBudelS6Yh9zH7t2+dad2GfzVqEFQ9vcF4CN0qhKi8ECUCAMSPKpvu
Iw6KioM2xQKgjiAxu7GOYEJHOHVOBWaQvpsALPNg5TUgPEJUHgBb59IEQNNg+ZG4UZm6qtzVS/9Y
KlovZFg7Z18svPiRT6KnmMiuiyRNOf81zi3K7ZFBq9o70QSz6JahIKr9OWnSKiRdLlPOT3P7zyQ3
b16I3FckV/OVERnOK7o/1RfEtvaekOerjKDRo3nALugfKX3YNg7okKJ2Rmmevx3HDA49dBrgxv6D
uSPWPs+IOKnOnVaBoZqtK7uOV20sngJzmuhUcAC6TcEKQO/MqDlP3IvUiAfac1ty4tt+sLi/bj5g
6z5GYgH6wxmuOeBRireHuy0+qUmybYMIweoUPP2LeO+lWE/jeFcR7dPUO3+7qdA6VXVrsmCjTQ0J
z+ZoU63z98wPpLqxCWgDCxzifbahrHZqpgKqwiUh7AD61YIBROejP1JotAc+2f6BtwXA6tdXClpd
sH0umkRqOmZ6Of89rXWhQvDX0wi8+aHRNKxLsNnGA4eXtfc+tKhypV0w8PV7MxVze/2qv28OvrK1
DIHujfESjElZfWxZbRMwlO9Au9IK0lsez2s+ugKAOBVYeHNhBt83vUpCRjjuUL98ksuR5KtLsHhu
6HCIJjg6UNMoNVAFznT0NDw/Bl4GwMgXt7oBtxgTqkYTl/dQ8D6oz9v/XL4uPPCCrBRPhsxaPNSa
4FyJzTziTT4jgPBBGm94wCn7zJ+mz5oeGjaw9x8iTBPSoHv7KEhUzpiV2INoDMLnNxRMMstpm7j7
BYltOILIgCobhHanA37fuj1zE8uNjwGMCUnqZ4owcfA/zksgKJ0NbbOe0gsb+aOwdDllffI5zfGZ
u29DI9zfcGK599VbX9VHAi+ePjqiFbk6/oIRUxC5VizFqQGmrrHQBUSyAPfPBUhgfHu1t4GeLWTs
s3r8m1FlSr1bkMX0WSdtYdZAC0EWlJupH9fUhviN+fGx7/KLiEp7VceS5e4E8REui4wgLtr2PojC
8Rzi3eenuVQ99y68+N3NSHYplCdZvhg4dkBjoIgNlVnrmGsbe0AXi7Yzyh2Xf/jPYzwGN0to0Fmt
93Adkz6cH0bB7Yxtib45DvOSl4tLgCXnjOcR+oaOoirX9ICoG3mMoclpt2DBUdH8PndwFtbjYfG1
qUDxER1kN6fubawG1VbgXzUZ11A5KFmW5W7GmTyEhq4ilR+67EUw49UYcWc5rqDaQE5iA2h2fzPy
Wcr7AwSwb4mBbuGmmsEuOEHN9OOVdq8ghTNfWs4ZASM/h3f/+IwRu2u6G7lCeTb9A/knK2wJ1F6x
IfM5MuONPwRFXTHIJJcJ+FB/IFmhJ23I5CYkJRcGnOCLc/VYYisP/cQ2dAJNPJc1feu58ahugpRW
wrpy9O/BWBwL/BaoOOzUsurcveI8MylhDHJzqhNW4+j8UmatT0n9YBFS0u7bFDX2jEa/GN98Obi5
zSqky5/TCTc6zs2/wn0Qx2rjdlAEjWDGIc4yvDueERT7G/ASpaRK9mz7dBMOtcV+Fuaj+/5cE83X
hvYYs4N4YHS9qW/399wd1cz/wbkgJ8IKK1W2chSk22i2nmN0gaNKFisBazX1OcYG+PRSUqUqvjhv
xgZoNS7EWcTkrVxzC7SNp/VxRcXaMXi1sDY/lhRDWnsKX0gU7zRTKe8ARfUkotasNIhKMhjkfiBY
sacZu5iUOeR8nE3xSIKS27C5JdBPFGKnhyQF9heSQq3Ghkx2ZYj/xNShE0xtwRDzNKRRsseau8iC
ZroLbriaEh9nSKsijjuXy1Xw2s6bnHcfHUYvi6p6PFLuWLY6qhVSuv0oHiz9Hg922PQiinj77SKH
NIotBLexCG7KJoKU1CPxGCLmbz/XLtHOHVgjNzTHven+Ycuw1BvbxH7a+bn3KvUZY1YNB7mA/5wq
O8zp3PJprtC9/fjvVtGTX+EyA983Q1COdMtJ8R7TpwGidZ2yq3zPP/cQwmksAYP/SArVkcvn2Gnk
7i7UxqQMv4ouEP20AD+o1tYreUPO30ZzTwvIWcAL4ZpjYhlKGOm2NvDZ4XXtXEYbd0mtOyVsVJ0M
YBsBQx9+dAH9fPjzDtzBDrJ+yABtr0dXQ/pzPJeohC/waQaN1I0V6hsh4pOJoDRcd0vfALATe8Wd
RYCTViNASoxTY3ff77XS3fMTiFVcoURm2ST484iFpiF2uACWgZzq0Ig24/bzo9Ki1oxnYHJlveYr
UE2VY1ci9FxsThJxJhTJZfAlrsTcpmk/WZ6tcSBiRLM+rBDZmD7/MGuUr/VkG/Oif1y2UJsak0f/
IS1hilBzCExNsORAJfmnGWXXBcx/oJnquJBg+xCIO77p2wNq55eLIALbO+5qpJdZ4TIXvHv/nqu6
YQGET7T865u00ycsnH4iv5oSPKcvOhW1JZiSXh1WgOIeOb9f+klKWhjAA8Uc4AZL8AXuiypauX2w
ViULpVeI1UB1O6LKlkBF7bs7+QpUJciF0Sj93ppXB8MeOzUIcyTzJAd3q5fR3YUxwxOHtgFbz6La
fliPGEuKPJtQKYcFgnIUiudowlGpMgizGuqAQJZXP15dCZd9PtbiCGGzDf0ux9xxpo3HF9aujiMl
56giOFXYvSTdtOy9yYC03YbXT+0wwgdmJ10CXZ+loeoNIqwWVRLbS+6r2ZZ+6wzTSt3M2N6SNT7f
zI195oCekh6SxbNfvsJf1ifWY+mOTnJQ7yZjjksbfTH/PY32pk0lBjribHo+6CFHMi/oVxE1NWx7
ighUSvedv9codn9XTL/+ek+dyXgBmpUf5wV3I2sy7ijKdLNv0jXNLjCjB5qR0PrZu9MiJMT+T4/1
kyYDcfvD3NfSan8lM79ryRveuQJcHgIK+lFi6rhbKogKQz7E38EzVC0GpMfU2pmzLk4oUdveu2CT
sajhxepCjaddyUiYPZhJ78ngNof81uPn5dp7d5ApBDjhfhZOPWczTcIyW9QRaIt7nF9+Ezpv52AY
zXG8dI+9Z2+lzJqjKQqLSIcsXfWo8QvP1d/EHv2s+DHydtK5WRVmr4C2VZINsZ9EHcRmVaR33bsZ
yC63UFPI1gLqQlVue0IXWl74LrQjka9wSes5D4ieVjfDGMQFvGCvj/NQJiqH/+myYBm6vxWeZthl
6JD3j2bIrgeJb+lx7w4IIWiMwmNJ177WMfNf5Io+PFhxPvB3kuhL5g6LuDas6/tVafoQ/KY2AKQq
fcd/TDbk92rbIzxQILHwwLjc5stWKAwsWw6rpcTues7jfuHGQIxjTTVVoo0kCdQ4BoX4jbaddVyp
tZ0DBRm1MnNsYgIODWwgw6d8WmmgzD63ghSLMPW0eTxy1H8+rbFfba6pJcYaT3W7jb6ihoBzgy6c
29mLHPRSRWP8H1vRd/MVLjcojQDdbTjyZgGhMg6mmhoRz54tNtbFR4kXRQXQpUCgCdGyhySnqEHD
osg3FUPqToXdIJw2jBWq/VZbUTk25UinZK/vsQVr8BslqSlWLP0BaEQZAIN4kekmB7ZWa3hMWb3J
bRYlalLjbmPzi+GTXI/l38ackEjAIDAUzPQDBXBLrWHk9GsT+i5H2E+Ez0loH2AXGk52XKCT3E+Q
IV6j8v/Yb68hpg6E9Aacv5HgFgnteY2HOQ6KqelOKE6qPkWPLlHIU6FFzYZdFRQXflZxFJQGfnHl
r7wpQXjZ9/zsq+3+DrYnzD2i7ssuTpW4qVQ5bf74mVmc89+m9onBANbLAynif45eAtdCPzaCKHX1
9M4pfMAskwdUtRCElbDOo/kyeLp+IKlCyUNIOBHePjvkX/0T7jhgAa9/+K9447v+huKomyprRYal
NscAcn0ZIxuLJntaa1KR1Lh0/MDzZy3AGw1cEDBZJ+FfQE20N+v/xc5W1SBqMpyKM+P9GZKyjXc5
SZOqBQWp01hg0tz6W5XaHTcch9XUA0mRMr7+TC299SwrHMstaB7AKG+B+RmxC32A5OaNASwYWThH
VxJY9qzscHCh7J6JvCpHr2S07YYngDiAxBgGI3epwr1R0YPRuA+Jyrunj7CzmvKtt8x8848PYpFB
9x+LIgda8r7PSMoa4kCw6vwV3qdG4U2E6u76+gedp56W+rXs0YTzOwypdwLpEYrxVdLMZR1cF+MT
LLaMlB5VZLn5YPQH68BTp3o46Mm1o2obzdLrkI6ivUG1tfJgHtDb/YMHxvyRCBLHnyDXSn5o2++O
iyHLgeMZgSLEp+DnvsJyFbPsCLyqorV9UyC8Dli4hmj8SJbITCijkZTqa4lXtsWHWDcjDC4eIY0U
tR64KLrlRe8qGZkA1C+2WWGQhPDkF11R+EBnJID6PO8Ly6NZ6coOLFjifNdBH1r7iM3D26gNfiRi
pY01iJ8EyZZfSuGBLdghiAwJj7JlSGR5IDbFKvtw6RIvs7YuXjec4VehdsDCsP2W2CyDk1zj3sEK
2jYL+fh60JDTcpYHiOJLxzw6VKKewEpgYFin/vlJ54mzjqHhDhCc/QH3FqYWLxJMBGw0I32kLt+l
weHMC0ScBzluwLhuwGu06xBEGbls2oqV/q0L0EolaD1pZZi7WO1KKWZhXoHylabYyaERuBJ4FU6O
jgPysLomYugG2HGDA/PeYHLCNvKnWlk4wRa+QQEg+iaQUT77B3xT4bvkTmkdSqtX09fKW6/AsuvX
QDSBW5gvsZgfSRbYwuuPCf55hwM3SzmLawk6ynRzEgVX6UV903UenGyGroJV9X8/Zh6rnzd7r4Xq
heUPh+G1l1c2bjHFN054PLsp+aXEeKFTepYNXXu/s0RivHhd8rMxSQn30ylfVHiN9c5zZ5TeSI12
a9ufVFljXfWXT4NXeA6p/kD21ZZh09ipagtgiU0xWTrTj+GMC06hsuzFvhp5E40L3jhCNfOWjIWs
u75Lzdy/wDGdBPeQKlCbr/4cNJUqzNgEG+66M6zQAxZQQySRWtQwjsEVdFsp+0xefmffIN5y1XNm
ukTR1OvjSNhqnhjsrWojz8j2JKuA+g65dBEfwWgNvdc6vxfSox+2eo6vnAayLtcP3KolSxUpijxo
AF0IGnaBUypJhczuItFUh6Zk0r+/HHvtuqA1ClhrQys86QQaNvIRP1Na6RGe+mZK2iDE0g5cNBce
j1p5pxrTiyx15SWEGknPG4GN5TpL3itokJqx9duDth6UfAwK/SV3D8iMK9x8F6/5LzizcMDIxs9N
H6OTtvJwrrkN1hqTa+j3DbRBJzf/5YoECNnGPB9kiS0PTLydfG/BrEI4kn71TF1fzu3g8SdlB+na
n0TnVbh6tMakyXnrRc07MmN2V/+UkapPkLFqPu/4GsY9oprhBzwWvEhiJlaEpE/nu9DRZ8iY5Ktj
77/VBmC/rqAIrrcGtOo94qHa/rhOlWHJx51kgHJ0Ea9n3IpQvemT4DQNpQqzW3exBNN76aOim40+
6POH2LQM6thulQ/RNNjuSHy3X3j8kxy2hB+VHdnNwwOHenfnnHd1OmpfvbYIakAXIsuxbyViAtK2
GywwZLtDIAn0orI2fCCYhQprwK0xFKVI4qPnx+5Bq0tQa5U2cqljzovv2cH4uA0Ujjp3abJJEW2w
ip/O6d6djRDCczeN9j9iQSwQ0ElqZ8MhYKCbQTJ0NMlf+V5yzF92BPc0Q3KztTwrVEIsB3vCWwo/
zNs8DHbhfpoVLdAtEmW86pRHSrG+xl2Tj8qf38JqK4RVt4okUsffcUa6er9IIIQExLI98EFzQBPA
DATYj09iwdfNhrGX0uVcorF0RXfzfjRh1kVp0cumBxppnd1UWbk5ncN5mSoF/D6ly++65t1KFVuc
jlOBDAgonhKyz60cso9O9ag8DhMJkfBIcPf5cT5zMhNCr5oW7ntHVf9y7CXHTomQwT83IbNXiOz1
RutyQ5fkPF8xzXg/oWVsr6KmWNLdJ31DIwmlCVMGxVh7fTmAb80sILqp/Ld9IZklzWdGth8W4SGq
3J+zb3lfSpxp3Dqm8qFoZ9OGvZMEVOdSgO8ZmGH+HsqevKQO5WUj/FtKzMEkKx4XdfFvP6U6Z7Uw
1kZf6ugWWoopu8Vrw56Nbj40ZpqlemJZsv1J0aAnp6/ch2KyJzA9firhdtw64OGfyguwYavy1LL7
VrbmIgJXjthFizYyy9sabnzNGbqgK9kYUVUhrJbxV7c4EY5fq1NYuwWJndhoj2J65nKxs9g3MJr2
fWJEh+QwS3UtRAwBtmXNKxrdrk9J7Wo6AOgj/32Y3NfqnDyqpIxs7BAglJqSueKuEGKE93em+lmY
qIguPLfLwQiBoTJvCy29iUBNXNVfP/1Lnj0Le1ngsAjpkT1geGLoqcxLc5qROcvkPF5KgNcnHTW0
MIZVu9IpuuhqQpBTE9gEA7HYfO8Lq4A8YUdGFAoJ1+uKBosqWybqea/IU2tY33sqCCJYG0J2zxcx
VbaFWaBZXKO0zGx7wRgwKLT8np28sHe5EBJHGIwMA/bHjdkzJeWfQhYT6cdpJDJrh+406k8xis+g
829DYlG0wv8/7mKPuL8CfI9XJJugGoMOVXLKbhjtnSi0clipofQwcTHMJaYBpp84ZHEJP69UDQvU
gpnckr7qodN+b79SvkBGYersXGKJlZIUoU4FGdrnPUGEN4vCpzK4kdU3yO0o35JFVShhyz34Vl8J
ug8iq8f4QdKgIs5SEaRnuxhr6mW04voipHSL+4v12A+TDcQtIVUCfODRjCOA2thYIkmd16X3GCB+
/Lu/pEfi1bY2lTunmJGjxIgchTlEeCADlE3t/jO9cu9AK++jK/mRZxYTx3fYttke7qgRZwfYfvWV
EBhIr+l5G+lLcLSY7FhHaA5piGV60zHCZm7WLH6dGiOjP2Ei8vGGgdnLvpqxGe8oQnA0xkpMR4xm
zjaUjAL5C7pCMQ99aXviYCrAFHH2BHhQuvqc+dX6U3CJIuMqRM0JZT7fvgzsJq02pFTGRwDO6vLZ
HhxWkAUPpxjc+V+aDNDQ53VbwtetA5VjXW5R5dy8paNioKRoeaJPypm28sp6HYKmt5N4jFDn/bE3
Fhj4xBKWi50zwgyoLnIJpBoxEOqr+7u5jnsYrJR0ziUS0/FtIOlocv0B7l1tqbURknoivEnVUmlN
L63StWKh2HeRZ59zGPAUoteDFsdNr2qkI6erl+nEl64CfM/M9/ORJM0rm/pjuk7TSkqWPBeRJ0k0
JugvDaTi5DnlruvoTI9t13AWmgLV2D/dWF84iFGm9O7+wcqoBDNtMzuqp+kG1hCchdVzOuDZAX8b
yPqaczmX6PMrfd0smkBZ6PvjuUUiSIL+oSDEiK3Kb+BO05bKoZm5CRwPTTr6QCKutpNU3yZ62XqB
SMI/LjdOeS26MiS9gucQDzv5B03v2zwj2hyi3hMaIv92KcPjleqCAAL+6YtbCfqEw7aMh8ZdUHOO
ROwcjHOg+eV+iAEzBX2CGoVvS5QGmCxy86fjJbGgEqIOMZlVWXz3w9FpDsEokeQOdXnUN17yPaJs
q1mojDRXhoLqEbhdBRUbUJdtZvy40OMu4/CrAsq19TTiEUv6HKaDzi9gYK39fkzOCio6W24u9Nok
tFL2gYCNpAmTMyAIJNf4IiXB+ZEc3vtHu4jACCLOsMW6dCIlLG+6eUxmZ+5pvPtYrO3gIwwzrHPh
ifV7VpGJ9OA9tjK+08qqa4uArrM6ViA/mwV019R4T93afZKzw/ZX0LUJWn6Tjo3SvHlOrCBfCtpC
bpBhG5GCDuAs5ulZVR8Z5l+BZEsCEgW2qS7B6fp7x/kydvzNb8GHiMepevdqzrWSeF5YYuPI+2wU
Az9VEENvU5UXD1fp9JtaMuBHPpSmrq55ux0E308bNl2hK8jvposmYJVLQBJDXH+GwUK09LJiad6K
TWS/pY1ESmXcOD4AC+TyFwsCaB5bnz0ezNLc0QxsvwVIm92fC5WLtgY8KVRdMIuNGhYSIqGsmINb
t2My4EBI6MWh1X3jUlyRJmsfybUP3nca7Ps8m9LxhPiNoR3H66zjwH0xvvtIFywvVRS7lMldXNFW
ZedWeGWFxf7qnRsJzxOsX8MeIv7lXiCEh3vfcJ6beFQwtd+GWDPbTa3/mFUobCwaCIT8ajzEGXVX
T+2dt1ZL+KK9Zg1igyMcyu1ghjG07PuZmX9VTia9Hopcq5yTb853ydSkIfI41cOrzQ1XQ4MM5Phg
s3w/KmNlgbCSdDWUggZ1+YPflEvCk2eHMixhHz7bnKCMICHvRWOlxUjQUdiIMLePA1dEkRe3j2bU
3Pt+HaoYlYtp8ZH5wTEm3g++7WmJTxiNjuxw/fvqN3C2DSBg4jZTofqQtEaTpi6JFxqCLR/o0hMY
f/9sFtUuogYDly/QwTYZ+8vl/bYe9larq6yNFn9QawkqdJv5cIchyf56MeQ2MExHN6Q3TBwBC6Ih
86QRkSpnJMDt+40NHiz/JJ4/N6qsRHYcd3w06MUaoITatDrq6zttuFEGrXhOTHgo3OVPgWGXbNeL
dAE/YcnOh/bEUNAJclAWCfai0aOAtUWVT/99otG5j/Ufd/32CRINNRZLNREVAjl/BRyza4XnobDv
LV03qyRb0aKA8Lzss7yI8SUETJjBF0yyqygXatgv/jZQfo4oWMLil5ARWJIM/qwOw2PczWgs6hvi
BJKl3uxvvbEbsQ1FYnJA5WsGjqRwcQ2gHlleL31DVRQXMVzFmgusAyFyK6ZpiRFEgM/l3gxposIq
jTAfOg6RIAMjCF4cePDfZgV/ZRY0hpQVMfC3xW5a2rh3ZOpPeqyMm+YvxbR5lltgIw6jTBsCOnxB
LLImUf2JyPodId56WIC4p/d8okjOAOJxdaRD7dT9Wl9+YkYeNZkhzn/S/h0pQ6zEQK8i5sMIEaRm
BPdSi2ivlIClWCKJu1cIve2YUnrZVrrv9uJyp1776Ta8CV1mLoLJnEi07vwsuFGPZPQf1zfsOYyz
+gFJqDWK1K/V49i+WH+YOtIDzlYbaIgCe755/kml4PhB9WlG7gytTU6nlXDIGEQ+SPPb5+k34Rns
Peiud1d7DKcoeuc8wXy850LvX5iPIsm7Nnz1wsHmUjeDFnVOSYcubs2fYj/3kblFkKUz9veUd4U4
SYsRPxMMFQuMKHysi0CFG+ojPXXqP5sSgV2D0B1orCYriQzeOeQjisHOja5pD2vsDWBrGc0/s3Nd
9qgDcSK1fT6Eox6ic+H8KBJxIiCv15XM76G71F/63XWLWHaZhf/Dc8syiSldxDf+IwAUX87MfpQC
EJKmYv+rpjLn4oeIzykbWHrAJ/LptqI48ho56vOVWWHapBKQRPW+6DIgdRP3NQREEB8+L7lI7tnf
+DuyGYib6BjebUef7I/BZK4rRuOdDDWYEViti6Ec/r5IrA6oGt5NkhQlnWdLw9fF+yyJwXyR2tre
baqeV0u4oMFW4dzU2iKX+nUwm/U4+7EpKFpDnR7aElBG2bzHp9eX/8kv8BsRlyDDrhPHg1EUmAhJ
Jr13liuuSr3z+CArK2uTxcepbdVeUtwO5twcAxOCfXPUkE1rQG7pVjrGCn5ynHyd08VdxtiTDddL
lRn/3JdCwtCpjb7jnE9VKpOVluNNm7U5ADem/K7YkP/rB4UeTFOolexzz4BrKKoMUGZc2vvvlGzg
sm9kkGoh0ena6dYXSRh6wJWGWyZd2dQtrvJ7+5TIpeJjRw0GY1KdZi0yTeukdbEWG4s7Ceft/NQS
nG00GG7oH+D+n4/Q9pMF+F4bmH0pA3b+KWN7CgFWphYaT7Ifxs4OTMAj0fIy7mDAm+quZtNsE2Mh
AX4zm+AqBtdN32y02oxaEnonAlGwsYGoJlo3UrGFSzrfeKGLNGk3geEZWXKrhQOyScqO2YNiriZr
8LRe+4GW/TNxjgXu6TA47xX/IEWXDYU1KF2qKvW0+mXW1PUVh72wt37hIaZ9dAVXiXpiFxeZtTql
8JCH8duFg0T371cRIHymO2hiZrarRNVzM2UvKkEJGC4GKn+DIWk9dDmLCcQeRPcftRCwwhNtHR6k
9VZDHOnD40nO9JBC73nakFOMkhr+Zylp+hqfT1vbsqdilbV1yupIvHid77TRzXi3+CXf0ghFUmH4
MfZjNGTbzvNQ6baFZImaR2Q9KeGrv20Golkvfzx+3h1K8LNgdmbCncZfFqGZuIL9OZsF5ttlQ3H6
STnEKcy+tu8fiPkERbnEk3+2XMFBbcUvVzLZ4obubLwtch3VKDwz9E6RXI8LRrdgd5JWWN+10DsI
Zq3Rg42cbE0Eu9NQ8kIhxumWagz0gn0oKLf25jqjBcgTT0LjZP+RuXdZDclXLosA2TI9Q4dIDalc
TZo5Wxa/YCNpkvepXq4rH37apUBCj1yO+KJz121zertZJRUSMwMhu8Z2s8FIuNe6X0hBGd+KfEUd
96IwRYpRDpAXaSdRtlcmAzkv5mWTJnTi8OSU/bG98U6GV4kwwAe+h3C8sZwrHcF5ioprJKUhoze5
Utd8ln0gdtxq7WWb0SRxgqBkHGYM4M182A8oMkW3rV4DP5WgYU7Z7c+YQHaBSLhQ+CqEnP8QkLQg
fNuzztgJPpYismoctQk6AOTI4bl3oaQq+lsGNObpRpdvLRmgb5F4UOty6/0N1Sq7h2t2cLicyjC1
JxKUD6pGTmp991nb5jTIbiKcJlhrNYEznAqxxf5TUszLC4TtUO5dIre8q4M6BEw+bGT4Pty2G9PQ
SEZwkRKK7oxjz2fl8gopTZjrD/1T8oc6t7et2bv8vnc66D2iA0j/fw3MxD9oR78bMmohWw5qxGhj
Xx9wuEjCuCKkWmhXvlu+i9lAzhOUriR2KFTZYaNuGqExugq8mnGAbbUyq6HAqmWxTYN2ls4h30cl
5VOx8MKOaCQ3x21FyMEBbrsNvKY4QDHZM2l7vPUavGDCXqzJdCqlIuEiJhzl5+EaMdgTITAy5dJN
gdbhgwlRhVWCiXtqTCx3s3dE8kdLQ9H801ohuCPi4ChXBUwakIo5Kryori80jO2HZZfnF9nAmM3i
LTKhLYTMfXig8ciEt3oUh0MDlaGQU9M1WGWqyOC2wzBKfN2F2ZAiCQlbbAunBHYFJWcANsicppke
SMYZYmUEBhmPlN2QdxT9GliHJM98yu17rOmwCq7Z93lb9bBuEwLxhKAor/KLl7vsExG5JHv3B9id
HvZAC9O4zwFFK3Ks5+G7COos8VFDM8G/KoohkZ22p3EDqXgW1I0TY1GyKQTPq6gNHUDYHzBpxLJ8
mGFnLQpBJYiOEffWslQXqBpjAgXG17qj6NNtKPGS6BM+cRKHSM5FndVFDeh1y4WVUCUenYPYHrZs
3ELU+W7Z4VNVMpfGnSBbeZwWUrfmLrGXHdJ7W5u4M7U1TvXE7HMnRy95WIdcRjFjz/90h1TB3GR3
hhlaRkShUz+hhmjUzQ/DM781JO+mqhauqcHiy2943A/VS0fyjF9X82R1hHJW9Z6PFBTcXb40aAug
+mvuiutIZo0cwjlmJHuPWhbg6HK9oBmAZhW1BaSUTf4NJXClRDvJVeVYydeMw7KsCtFl89pJDO+K
R/34khoSMwCmkc9kXi0TTAU7PRvgcugRuYVu5BZYwA0coUL7zhLPIijNaIZ6UhnBiF6gLM7YKTd3
QN+VC80ZYZ9g0P0PungXQc+PkdxhSHZiSy9cxhFLIT5YeQGGjHVTVAaQwO3ht3OLw8l5dZqceNom
/wFlEbKqON6AH8E6qW6MIH6+p8BQTHdcwpU3U1+uJaRrxLO5hvIiJsMvlCP8qyZ2ZlNdeeyazTcM
TaXcqQ5SC2wpk0oskH7HCwBiubuYpx2nKEBtaYnx+WwUwJHTIpfE5aMgDSlttyr4a/9EqbY9EHYh
fkn4aRtYHo/fuVnCj5WYowTs9vfVfBpzqT9xPAcQ+anGyJvX/iDgz5fGz+ohsi/879RMoW9LYHWx
aZyanKXRgdh11knP8DIvxG6zg/DZKPKyFGjFbcCePPnEc3poW9bM/tRU9BOMTZl6mcVvafQdGAkd
MwpQ5PnoUj6S3Acg7s6wC0S+jY4y87OXwQ4zrvUmMB2Lc7neOZekRLWJnEtwlRjQp90sXEPuKJJD
93IxHoQCKlKlIPlbozucxgTxpJXjwgLBijsQT+wa5XzV/FrbQUQvGRjLOnmgd+ySHTdj4lYCdAyR
ntv0V9NrdnTtihn+7qi7FJyTNNzGfXVMNmrgASJ+x3lDu76mUECHhtPg75ggvpzhgKlNUJ2Ocjdo
HV54JNgw/HX/SmFsSnUmr90a43alc5B/bzk1tYIegtAfwr2dy3n7RrVdrhC8QMjqH5eRPHjzikWQ
OiqtslpZK9Fg1MOdiOmZRxcg035N9UgkHo1TUYQZ8w/GukqAW6n8iMURN9DizTKLIxX5ry5ulxtk
mLFY/THYWDapeoLSbC2q2+IJLb0c1DmulGSaqybGDqv1tN9sMOZcEUfxWdd3CPXSFMXTyrDyzO1C
96dnG++/Co4K86wB8CwS+ijhhTeXMMNKNxL7NSls4s3ZWX6O4gEXhCB3spSTvkbuj4T/4VFNLhdk
oPluYSvp5i0J7ZYJHFLjsQK3rtUnwi3WiQA7q3zq762yHPeLfqseFXsX89Jlytl+56uLelikIXsr
OFGQNg7es2x9ohejERhpoJYlPR2rPnIonyOA5Ngg4R4muHH1dQkTpVme9AScjyqwzcJ1iBsylIdk
TrNkduwLWKRzPpWKosKgxM3Df97JnzJpFa+tnq/TIY+vApnpaydZFTq/ZdKlQBsWk570Qyjho0wy
pf/frmUZcl0UZQTgekJoiawa0QOOThYHh1FUb4ddHWJBBZcQQ4eKf4+R/4eBOa2Po/nrxBSBg1Re
N49JLsSxA3bDQd0H3wSNDpWI3beSux135+2ANxjeEVs3eXddyAmoS9kV1r+ppLsiijg+h/kpffkE
6YXKkrgYa7lIyVVu+DCKmZ246XjDxExqpMYFP86sJRLIRZbBQy+a0hBh04I60B1vld17vPwkG1Vd
N3FiwdDe7RD+XHjcGbPl8jynA/Q+yPVLh50Kt2fUpsk4zqjfkfBQarnhds401lXwfWEcPvGbnKln
qRkO7RuJhyV8pqM0qZjZLwG+htW/q8CDfYVJ88un2L+rzyvZPD7cWuV7sb38scAYIUXwt4RXWsjX
Tp7bD3b1Nm3pR9qgr0mbw29GoOWX1J0IjnbSJK353hHYZiKzGF+EZK60GudcKKt7zeyx2WI5Wxh9
5RcSEb32dUo6ZkIEIcGUzpss4myszZtxc1QbAWfFNiSbepdsISltW9OVqZTyltA7g1BocMVsUV9/
t1WwbB7iYypqTo3oRWkGnJcIdGisDO5UR2thBJgRqKio4pi3XxH32OQtMERMRdva5/OUI/tuti2F
SSX06DIacH60sc88oyztXtrBxCib4SY4e0r7S/EuWol4+uyIFGUe7ZcrLQ4jQFQn9TKPq2YlVbwF
If/zWnj5pm0fY1YEjfCLWyxhOIR2BGEmpsBNWNqH+Ah8KOngLXmir4K2Xdqgu1CkobfzsBttp7TA
xQzHMelMqNFalk82nPQx9zA1QF1QAsY9e+CNzSzRQimWZzj9KoffLUiY90zA3tBYtAO4ziMv/vYT
9JK3B5ex6w7D8sfYWZxFEYAYWfP3y21//ilouq7TxIAwXPSzXF086w1ZsGivvGu6eeqp+rMQib/Z
NCu6y3Z5bs5bgeSpFHwC84Z2hRvd8gLo5qtUYXV2pt6dzp3ohO7hkH0fyPE858BE60LGZ6UXnnTX
cz1n43Imhn4I1dnLdGj10RRrXsEx5nDQA6zgTdpn9jXxEuIIcrZ3kubJaF4UDcu+iqXg/OtQThbi
/jQtmdyUD4K2DutoHC5bUUFnPPy3jXk8faTzTze8CA3en8QfLeKwUZOOlOsIutBXldd+i0iXoNez
szppvTIyJUQo39BoAO6KkrJmhWVVQeO+Ye+NTMUnZn1SN672tIBKQeaCSMoPIxFgpC0IzYEqI/bA
FmaLqs9+63YMQ712h0M11//lgEH6xFQ6TOsUu14qh5z/Gggs9AQfUyPjTk+Ss/jtiAuzBFM5Zh7B
lwNIrL/O+pU0Ef7zZgL5Vqgr6PVfSdAa9hChGgIzrWFiBLWyP3tYW4ed/a9VG6eArGWldsEDok9m
QZ6gJmHTZNBWsmqaeAAjTZ0ZNLuL55E2k8YFADPoFbOA1q6SOu7/F0/qup981EVEExCaAqzbQ3Fz
ICjgcNM5LnfBHpQSqENVItcd74kB6WBoJzO1Ij2x9yUHurv6M6og3dI9r37TE5+vKmrDfzCxREzv
3OJ5pjYrvEBdN1rekpmQmmICQAmKkDQnMVkX9nqQ7S2j0CQ1bLCFdUi2CGT2CejQEfcNUC8UqVZQ
knSeBvoO7l4OQAf63EzkvNGqtwv3y5W2TjETqqDXDGa+Xcq4sbrmFrz8IW/+mKwkC5pnqhevM9Mz
vI/5KppDapftzCxoRyYTtf8OL2TrlAhQx3ATSRqDOdzejYTOwHNrnvv3npB/evb7w+Sr+FrQhiu9
4NkCglKAW/yA/7Ro+btmEYf+0I4Ah/IxNQfna3W8v7jJisnPC2T8wYnDUYiV2u+rYiI4Zx2LjaII
4X6bT4gm503Ky+gr84sqQCvNpLyXEz6INXTAV25kIZPSE3W3MR73v1Y/53PQLOdbv/5zYkGK1kBh
RjbJ5tezEyZKuvIn+XKNC2USnqgnfpQwzUzTyH1IqCRNIf2B+POOJKK4h9dvBlRlAQ3FTLtkLEt2
QBMhb2P7CwDqpGckliBHgL0ctdETRTFOrGnsYNCV1+fwNtxEb6xpmmFH/D1IT/2EjjXA5mpUxofh
u8MlRgGD1voxc/IozcEc0pryJgkhxAOHszldsN+8MGPpPA4K6AYB2UG8T2FKPRWtyCNtFb1gbOUF
+0HzydBRCIh6GA03FQf/vhwK4ZZ8XS8y8KUHG41VLzi20NnKz/dppl45yvF6RDuh3IFLfSd2fmVC
Z9wODO8A/Vjv3yg/kOSvYUmdj6qksrXYuBDY7vsA/zFDsUer+x4LUpHv5Lv7pdLPHm7W7mseAM+z
hoFlheGgqH9cohhgLeAFa7n9/1Niz8f/q2GfOzX2EIKjVecyoK3NdoCveGtx8ft7sPrHR2odt3LR
CPqRaBfN58Sb2dCIjUrMoyQhbOWmr7CHMt6zVSoh6STqJAw8KWscy8Tk+pyclx8zvhog8afGOdxt
c0ZRuanbjo1ObM2f5PRCDqGgDvkIcGxhDUh0dAGz57t5neHgdHeITpb+yMmo+6zcjXagkNeRZiPs
UIyvRPJ2yQJUwjbBgsJNCa2/6Q2IXj3egC5+uyarNCaKevbfFYceBlQLa8L+GT66kO51geqMYCkE
o3eEJXvTjn+X+2XdzjpnbVft3zWWGuCgvCTplLh04Ru50f4pxr8DA/xrvUst70K1fKHVhjbkriip
B2JfF5rSpfpXhCMxq4rVAT81wdqeZcN2bZRzm+ra+hJq6yIKTtKMJcC2GqDWloe4at7+LYoZQ8m7
eTeZ9Ym6BgGMxDCA/0xOmgClwku/pqKfkHOCmM7If9A+UNX/JPqWxbabMFvBDemoXKdxb8E3AOjD
tV+lo7t2Y0jhKF8XU1TdDGYFzzarjTVQXkbmWTN5tHMYEsPMqL9KX3O0/TsByhIQuirPslNoHZlL
4WscfPV8PeTYcZL9BG2Wayl2pnQizP8wg0eOuG2oJTwLVbhOJir7BBnis/UsA3bm/UNMjlpIPpDy
9gKFiO7PvTwyVnVJfGOqRBux+vQJJq62c+5QUuINDcQzVherWqHR/RPy0l2obDnkizMhNqqVJY/y
RELQuETPBKKshFb6PEBHIGzas+ZectTyZ1yRDi4PdvggP+CmwHwXvNqTduuRGCvgfo5Rako/g6j/
WuyoIygCTaaTfOMlZ6VXZDa1jWc/ngvz7HR3+52MkXLENS0dcFcw/Ode8GF3QJcjliMsHoQanACM
YPUHbHMYRyw3hPX+wFEe5kkfyqlj5/gJsleSaYw2Clbl79EqF8mWJBPF/11teQAI0rJtuAgkfRXX
iCaTzRkplxV1UqdNG5FI4jjg1b3wzGpf4JTUuiQAQKLcPFKjuAZKT2jpEYCme8D+9IBcV2D6PMVV
+LHvlyfc0p0+Kg5bgAtwSbSN5kZeTPgN3c6E2AJDWibC+1LDwyDl6WBBLGO0GzKQPIw/fyfIl6Tl
kVx0GiCuhMUl+6mUGCAPXi5gfho6kABr8ylkVahiWh+tak3waqT3Ci4NlkdAonRiYYDURpL9CsDM
xCZnMyDmuBpdYPz2vJY+d/AqOBZQYtDJIaPeVvhi0YwuaxonCGQFFQkuXu2BVB2vJVxqQ61Gm0xT
AP45+7/ddFNnXakTw2rO3HhsL7NhgQmmBnnn3eFUwC2AhfVR/4vW0Cvy+I2odKirciLKJKNpxwhh
c+W7hjOHVc+RPcqH80gTDffKjmtRA7Tapoq6mp10wM0VyH7pBxGy2HhmXR6ahWbX03YQ23QeNCHN
7cAYJERKRhWUZBOafLDKCDRDKUKWx4rSX+OGDE+l6rHqpGx0Ngtlko8WYIZXGTOLAAnAyHOAzKup
GtvoIyy5ZRaKPGayWs9nRx2EdvsMj+4UQ3kUdMq3E8sDI6lzOr2bA928d31VK0AJF/rG6JKZO5Et
OJwhPajta85NB+C32j0WnEFA+GOv07vg7FuTIEEe+7h6LFcYEEOZr5xHB747YqeQDsGkY5kStNOV
Kqu4BV8LaFnj2Vd7zbQ3QPjraDvWRc9LE188gdj7X1cAXYkzNVQwsI06nEph/21jTfcVrEC8iH4Y
RbG5b3ZtNgqcTocKoKK9YQr6kHRk9pd0prq9GEzsDPH68qElwBHcEZ1IDZoPsM1fYklGf/r6SDL2
mdkaIm1G7Od3qRsY61H0IReJF5VYg5aChw/CuW0PoBl/tgrAwaca7BFq+P/+5hqBu2ZUWBUwyeRh
wRp/hguUGlGisY9jz3Qn/wJDg/bz2HvCqPDD2eifDZjZAcdtEXzC8ztfgDeMjcPvHWGsMsqd72nI
kFs1rjf4lV8DqGM1HdrdffhTHAXOLT3NQZGOwxfonRn7ZWysfqgDSolBLvDji/JMCvPBr2g/zICE
nCz4DXB38XABbVai60CBHnDLLhLC8G38iuzbTfbavOP/fGgWQjjyui9adkHnAobl4EdAVdoUwPyX
FXh2nE1tE2/svAqTDTGqgfPoyugpewAA4RQj6/ZUGS418CgekgK1TfH4VZlq3Df6iK/0GLpiApa6
16/vIJYshAcOGQNQR2hU/jZtTpmPR2zEWAJSa5zmm627/n/TRkZ3q97z5/5k6eYuxz4JHGzTqmlC
a7/bDG2ohbGEEtT6dIVLuu1bt9QnMSXeshMe4D/VdOK6bfcF96W0yDV+CtPkpN6r5U1ov6S222em
gCXZalHQ0Rd1GjZg3L4Z/ZfKCRwvzQXYNtORVY7KDr31MXUDFhZUML5evXMmq7g9UdLXrDaw1OE3
6phIvFTYNcwWHygcbRP2LbXs8Ujb1GCfLk1/gK6LrUvSdaf5nlRr9rqerbi5JMXC4JNyTNa9RW2z
oFmf8khZdHUJyUtrguGD55GnXLic783T2km/MYJ2zqx3N0n/MWx9tbcDaBROeoocX6oGmOmQMVGx
9CWroeOvVtKTAwS9iBQ3EeDHdHEBqV/ijhCmMhwupC0cF+rs1LLhC0wMoOrhVmKDCSitjfP/Ixdz
pTPZh21Sk1LIkyqmTWrs+T4AF1fa9z56xeicg40nx1jXzMHQeiR5rkD1L7eV1GJ3L6payUJbHIZh
fCXCg0IQ5l7X0SM1YSPmYTQp67JPkF0/VB7/Jr27dJ8eTHcevGkSkYFDSOMmeGqY1e1Z6sTYQGjV
wk+VcJuRA8DV5RfhHxc4diKqUYzJ87Zc+tNIbgCJuQifth3m4Hag8a6HuwXNxAXN19WiWZbjzNQ8
HwBigm7QfAVWvDz2O4M/VHn/wMSEmQD1Qg2jtyBuxxmH403QNYWMBliGw8HOTSEW9HqhKStk3O8Y
6zkMRL2mL1r6dhFjurN1JGmV/+zAcAwpr/ujddv6WxsvXjVIL/RGDFeWgvzu+jXSG1vwBIEliwkC
VYCstD+E8JFEUC0rf9jw38zqBW5foZTyuProax/6EwC3Y8ZJbmLLPZklw7KXUKVE3vn0+1EOql+0
DrP/4px//8KMb9T8kguM2mZpZQS4AYADT9lk04uzhIjD4nf3idEqond8VKlcH/t+S+ItmJ+A4XGN
sXdKOZcYK1hzZA67iIzocsE1dod4mCcXx6CytPGkuZnLl4pR2tv+NT8AcnAqp0fh5wMI+9stWzQl
a3Oc0+6ky5xARg33eI0s5uTgak7ylUgvsQxNaW911Wg2J1Mr5XYbW60PQ78x2TiaIYfTu47gmHae
8xCSokJtH0dKXbz74zoMSA8x2Bz3+5ev6kAsWy2vhUdauRQt2Agqo1pCFIt39oZvy9lN36dyOUKi
ozUNMEKZLwd3UM1dlUGP0657bqACSjDWUduLisaZ4dl6mz7dckBydBW5kQ+X9CmF6jBLK2pQDYxN
Mp0eWLhvtg2X2Mb7vT2D/vq61hMU/rA2H7XJLPXrl0GrKsIM93A/EVsfankwI2P4qcnLglevlQ71
o4N1qUCWr9V+7CXWDAgsCIDZoTyF8K+LhIIbdbT+maxVaGJv+uxhsBgv1KhABl56Gbq0obxQKt3o
OmDbdwr1d+7//YE24gO8cElQJY0rcIQLY/RPp7ZHPt5T+y8TFgChKC/eWQge1AykmS9VZLOEmRdQ
U8Et5yOr11V/aUvaZwfxwGE3edrr4gAzYDeL03Ex2F3S3m1drD7iM+k+JBIbCLa/t3eUFKvjhfOp
bQvEmBepBl8IK4zlu5jPoitO9Wb7cZfex9jZxNHaeYvLN/h0wEYqBJAmZ0S22GkB4yHJqL/IZ+u+
zKI0I94bWyTVP9b0Ay/Z5dczp9my7So11H36ff16oCYZhxpOgleJdR0J1JgeiJp+LdLqPo5QbXG7
EUMad98HgOp0cDEM7HKuV7YaRRwU4IM1jdLl8GkEFdoE9JqM20ZMn111+x4G30Pa742+vIqXkNZ3
+GfNEoyeX/0a6UV0432IMNKovaP57BtGD0GNqhfSoZ8d4dC0soKy16zxtyXMxxojNLEoOJ4td/Ah
hoe47hc5RkkK5Cj6dUGaIVOIbyPRzLlEMKHsci8Am9khkecv44TW4MKD3eRCoNkm1OwHDi5S+V8/
+kXgfZn+GlnzLf2IhPQkvuuYVks1LNxtQ9C4Qf2VNlxKdlhgQ09RDHu2MfFeHzo+rfonzctY+Mfz
rgezNUPlmDHPLlJYXH0ziBrRRhGd+dQ/NX7TXKnjCvfmStgFkoD3cwa9qTEHEYgGqw+MWJPiSGQi
gSUt/BZQxbNyf7VO4BCTzNxar6s2TsJ4YDkCRPw9bPQ9IsLVqa5+LSWywQGlLwIolYLo/v3ouSo5
WcqxDPK3QZn9kyDxL5U91afxAOVeihV/P3l10CrqE60sEpGI78Lex90Hpd8N3S4ph9sw+UysT1mv
tXri4VEihEYJ39p2FVOTGnC3HTQKOmVGOuobJ2dEpxm4ZW0yBeeHCHcfuSAVbZEMeNL5Nm0nSOhW
DCcoIthuJnXMEYaS3OCAEyReCOc4Ez0jwMHafQAN3HxRRLhCUhcMGWmQ7yJV1kiAglv/U0r7HOKn
rlkO63mPjHl1/JqlS2W81N4of5SmtZv4jds7nz47lavl3n4O0BqA50LgMiBarkuJ6hO8r1kITcuc
qTwhyEYqS6NUfnP/MNLtFz/zWeS6uwccVoSa+h2Rfu3TBn8mlRI0WG8BiDmgAcBp9oKWLmA2U/Wm
osliISiS3JwtymvdgCIvwGNnbAPmlc5FMcOrU08F73FChDnNE9Yy14u2s2EFQB1gHxVE9UJ5+8A0
6bWLCjlbT4D7Bq7OJD+v6/aHwnOoy0U5eHxe2Hlc7FJ1sJsh/PiZlT0jLhhRBFxJEpKnodJ0JjVL
Fia+eNTo53TJrD8X0a5Tl5NcupZxbAIktlRnwbFRkDc5r7CSc+bGdvW3HdbbUO+BKUdnRk9fitAz
3eM6qbMMYxUxqQDtGvB/UQkEGA8TkZkGz8cSxjVonD2fHTS3KaxxIXcx0DOP4M6d+RVkRlDFkBfN
ET6o9bvZ2+smBmfTyYVpH/7pe6LqUF/zWMb/QMlMe+em01POpiIUDnGTCRy5D0em967Chj/5X8QN
K9LF7QkXSDnJopk7MzuENkTRZhrIABQGoJBmVp+H2q+CAoU4QYkoieMNCTA49UhIWnzumtHIiV+l
59WfxNPtAwrs6Laf3mMDATFh41IVYef3XDnIWKjQL1o0hDeV0E+4IQhmcSryl7cog28sw967bB4Z
J8VPqTM2dWlOaQDgr55csiNHysDuEvgRUEU+XN2N/EWm8x49W2xzB2qUS1hSHAqnkbHek18Nc7rc
49gFw3uqtOWX4U1N7xk3hcAKV3NdiBgH2ZwxUl6JBPdZdCUdIGXuKJl8M/pNYUr1aw0BsEXY7is7
D7ZiBWGjZAcfjIiE9yLXpjZC/0yu6rLpM3BsjCocB/RTiKOhchrarR6r93QS5cN8NpaEL9O/CkfE
ZXPt/mVxDMwA11YdLrISzo799210ZATnHplxEZhGLt8O6UaIs+LH1xBwsk+n6E3FdpszBgk7MZgC
59XI1ZkyiGmbFRILOMl0VSwvHy3guY8aXGc6Eeh0p/ldfu/MXtQZc6jBMl7PWMUU/BZ5bnzvrLUz
ml8Q87dkHojhd8y07+nKJQQU3RzYivQqCCaaIix5oiSwedNcchDqmM+HnrCxjVKcHwEXN5hJ9JKl
T/5irUv/psYKlveN2v81Dskxb519MJCXbNCCqrwpg8pKu9oHr/g7ZnNSaH7e5ddt74F+tLALrUoL
xUupYOJm3Kl4vDYj4O1Z2aH4nigtX5F5KDruy8dSoDgEFQI9hs3hIQbxmJDSGZIPshzaklbxrMLy
7tq25Qlq+t9StgLwKXYhXBE8N8cS7XYBIDHQHghX4IYXixo97+CNMBG1Elo1KHsqmjw0GrMqWgb4
d8GYLPt1q17TbhomvhcW0+ZhXoSPeG/L4BldaEpaI7zbgiUxxzS+2PWECBgfoGkf7N8UoXnRZpiY
Dgc0yhf1yKl9zXuhOmpk+YkdgFWhFeryiqp2K/IKvgveOlOw/zkpnUfEYNvhDhLKV5hw6Kn2tpdV
aJdCmmIb8nu6fT+6awudtPayNcLe2SUgsl/AH+/dB8iZ7LP/XSqRmtUVIkKXgNbHuKVaLACm9v9m
6P+fOJjkJctiZEtwGu44lsQDeLsyyq23jFAdeTdkYxWLCQCT6/lhqFLOSrPcrEwqLIjRMmTjlN61
hBlfJewNzbrd/tqnkLX2vdU1qGx8E0T5gfIircCBYHoa1MTdqrDNR9cBmSeTsn7F+Ij7xIO/fIKq
uPP7FjwPXFp/8Rqzi3rsU5B/evoRwcDqWnBHNUnxsLhexQi7ogTUFAXs4fdUlGdR2w5m7uuF9OUv
lSLr4OJ/VGbXGIcclBuhm32rRsJ13xmtD0iQgZ8udnXq8JioG3IeXaLsjDVWZuvBKAeWo14bBzjQ
RJxdlizHA6cH03tEvUf6pXndP5KkEcG9nHSTVdnSQajX3H6WFqEYD3GKhO0KWJdj1UdoX2U53D4y
sv+8/257vpXVPs9qLZadzlx6jkqHT4PA76SmBcJ+Js2sQNlk4rLU1gpo283U+T1nsS8mlMcha9BZ
smPvVZ8otIZBILpWJ75JjhbJhsJoXQ0iYHl2xdkA9GVYwX2CAauHpzGu95mlFDc5jovz5w6wFNTO
josEtAf+BcEJjSq5IXzkLuaM1N4+aD7qKU4Yjq2F5tQ8a4fIPUMU8QqKjmj6ueB/DpTFckPGrXXK
sUKoDEfEWiJMGoeRKzLwzgL9yhM2QUqHeOGu5670CFeFxO532VuassjCpdC6SNQ3gbP2acAU+iNz
DrEx/N6OXW2GdxDINltlDpqmIHCgWHeyiy97tFY9VNZfOFUrKsb5AcYTfnehQqB+wAfBIQ7aWLwk
wgwcu6z/+t3mEwWIhvWWpQv5t86zQCg3aozrzKuPzlQjNBXHhtgXLCpAI39UQg88O38JFi4VQxI9
kTwMEnJJkWbZCrTTJ1o9HdeI4PUu4sQ2zhytOc3jCzTJDTE5b/VDslqHF/sO8GwhgIDBlh9Gsi4I
QvzdtJbeZNyJkrbyvVE0ZBm5Is6NoUtiONiEoANRc7PomC9W2Ni3Og6ZUWriRXl8uGD1Qzc8dGcT
ovcc+a2wPAHOYiBtKGwYiE++viA0ZD9ZX9nz547KjOQkoTfszTSECtBL9ZTSXHjhg/yBwM4qlVBK
ox/2h6IWY38sO51eYvQm6zz5FNmoYpROIyE0xwuzg53HvSE0NdALNiJ9ZZS3yRWI0mkym/saAKGW
Z+ZroqmgdkcxS/X5JnuGC961h2S/U/AY0IPT4b2XwXqKIDVm3+NbzQabCY5L3RcTFuZ2CBGzt0ii
K6lG2G2mb0xHJ3DAEh+3zxutiiLRmL6ZDCymjBChef1qdrLlgRhezcH71X9T1mdoi/wb4MSyOY8I
2boGEutjkyOHyS/9uIkejpYKyBZAy4HxuaQR7PqNHQ4Y11sVnp5vVmv9wsZl/08CRjHL1WH+3HcY
9L2nfZ+GYq6uK4Jgm9WYowtm+qYDP1aedOiMIPxKbd56WqrhgCCHEcCFdJSKJ04H+M3AFLGSmN6j
/yO/P5LOVg5hfh/GdryXXuz2xerrO6FQJ2VEbgBaUfCTib0cEEXJR/vB55gTPkHi4VAmz35nwGr+
2eT6LsMHWG66CbDesZJ1GOGGORs4nxHxZlJRyLtU9MTF0UqqdROhFueetJX7iGLFLdTZd7Rqvo0K
XDM7xxVD8rODEhOSVRfN57W/ohmfOdHSR3EPgtJjxNRh4VBK9+HGFoM54sEJ8fV0UbPZCFgkcMK8
j9pFeN8NgjzAtC2az7vaF0rG8FUJwREWSDUKrRl40NSCh+1inT0NkT8eeUs5WvQPWa70/Olgk6oI
JVsIMDo0aJ/ZQiuiqrcGHPlh3tJZrdjV+bFvurq2+vC/jpYzzvApeeNOHbA2DLdo3AOn+BEDDoSi
nOpGFIvNoUoGQ5ksU8S4n8SoCAlVDVx6ipFQ6zMpN/u3BzIIBlwX80h9zf7KOq2jh/FvwGkSngga
A4ifwaKtVToo6fNrKFa3aRV4asyFbRvyXXvR14aA4GAhN4eD5QuXhR8YTOVJYFVJG7iziGgzBfMl
bFyJgA4DPBgcjkJaghDn2DtsdcWSPmVYrFNkn81Oz8Wh6502dCloRM5reYK4gRT5Ubv86Rb5C5+z
TNDEY+xwqpOEt8jgZ+h5AuuuvQUTfoYabskACSvuFlsjI40diXGxQP6pPGNGatg2bCH3PK4utkmu
e969riSayYiHcr9+m5dFyvaH8GOmdqH4Ga0Ihm39ed5dK7LU/40Af3++X6R9C3tATqfSJGo1RJaf
PGDGeBg/mXTG6g3gj+8n0IbFXP1wptgoGZUdgrhlnbBIVMPXM044CncjN6gEQ6cauqcutfI8Js5D
nKW9V1ff7K6rDRO4x9xPauZwg3rDyfJ1BwsBMsAZSYzMq22ofnC/eO1FiuBdSuHgW6/3ghRNlpws
bnyQyhFMAe0pgaVeg8V4Iji3cGdgpYzEYJLKTZjS3lxIMd8XsgNRpXKcwXbrS6eo5r+QT+Y7cSJ9
C5/cHhmNppUcUPqtpFDL8fnyHIyErmgIqFcFbM2WCXDZ1voAvbUhBh80s59RYKS2szWcW0rqG/DN
H1DoQZHKhFhBHEXau5/CF8m+e05s+sDCLDh/lB0eZGmvofJh8KCrqX5OyG/5F1UPVSaBR4cmoCpx
j4LRyVcvAtfXjyLm8wDSA772J4APUKU2TrwNMKN0P0uwpZ37MmOd9O7m9hcmSpJfzmMdWN4UdW0U
jrdxrWhzC0ba9iSdhjH3eKCEwJg915PF5lA3EpPaB5t4pzjrwbDbyNUajSqsaQR/v6vpQ9EdlD/T
okKtNscQxLBSOD4Bpf0xlKvUvmoByf9D/blcOYS3MDVOXVZ+Qz9VxaEnxDjW8ofEQ/FpH6cjDg5o
f+e+GPBd3tp7GnY4ijn8hnwQOoGvqKwLDA1GVQY6ipcIBm4P5+P9AnlJm/SMv2UwmAtkoF8qEnYm
NfdHAvJtfd+q+t6IWKy9hOQ5Zmo+uX2IsGJ+MftYU7G4P/qSyrTqgB8BW5L0yeqamLrXXtgXCXn5
+igosURrfjrMG8O7onk9XdukKdZU0RYz47Bi3JGuG+T6ckNbaQ3nMGntnlLTVuIeLFWHBWSCNaTR
SvuGbScVN75PFcoFyui+zNN64Pjzb8LhbLsnleo8/X1mEQIbglNwKEbLfP+mZRN65maR3cEqAUcn
n1CqAsVb7CJZOBcDimX8gVa9bzGWdmcUiXqkJ1CAjB81E4XPKx43W+XZsmsGHTrCsW5taeXJ3xLv
wil5ypkL/sF7FBI5iqXNPS4vfgt+biXHXYfJSR8qm1HUlD6fANoY7W3Q/XqHJUuJx6zvVBhgh71A
s9Kc6tRWOjFm/emV2I07UvypIe1gntgVJzvsm2LbJyTGbZBXF/bMW6Cf8kQ82eoW1a/MM0JoAkAh
wII4igbvwEyG/pex403jmB/JNLvuMsAmxtpb6fv+/QZgMCHoj/1KiWj7UQyt5xzHBTPvxXh8ypLu
x5qjZvCCZmnLIF/iRojHBtw/4B33F/vEI5W1IiSGLLuJiAwJQ81Y7dm4Dy0wBe8LkiMH3YcMbcte
ZWSYhrPL2PkjCB7DBlsLK9gpzGE00axu6Qtz1hYWzSqSjBV7k6Vg43UpofIoc/HXBU7aAolwQF23
gm8OCPoSavxyK8A2ILRg909WWD5IYfeFwVJN+A2xuEnx1vAOQfIuBUvrOZHRr16dYE5/AM+kk/7d
JVPX5XKSCN7oQ6Sr2TtS3bxVr5hcRcZ7/vmUf7/olk/euRvdPC/V6eol1inqJ6iprnXwPmYHy8Yr
09lFmD6p8/hkon6R2QnEgh4M/BGmIc0TiEeEkG9wqFkgJP1x+UE+b46SHNQ4zFF1UgopBxbrJjzG
6d3W8rt2wdCqzmbTHcXkexy4y4GjJ9h9tarSziy3yeAYN2Sea1L1cIF6yunZw0Js+pXGgvqQNlMX
VMnVRFt4DJJt98JQGQMM4L1WiUbny7ZL/9FnhRIBjH4qK1lNge+9GARhfPlQBzZ1b73POFgAdFgu
qnUIHWZG2Uk08bvvPa4t2TKnipsfeDe8zouwlN0353lAe7bHI2k+duK6vE47XXLI5uWrNcIqOU6t
U35IM6oJE0Lno9U3X8bbZQQFTa+UJDaVUZBiGDrhm3cWCuwVIy7YHfU8slHUKpOHlWr8jQi3YNXF
4EHgOG+Jg2JkYABSEoj2ddqTqruj1kGYQk2QuQqkWrC+yaVNpzIzHatELuQGG5uMYUA/KR/CXdIp
VV9UKS1SzjmLN8yFvn1r+Nk/6YfAnXd03Fkr7PypuxYeQ3CHhIQdYev98kYnzt5GnFA3fwqJNJBY
JYqxZPl5mNXHkCyp11rVF3VScbNDyrXo4LxKMU3jaQ/1nhcKwjvNaFCPT00v15Yoq6WiJD+cMikG
CHHWC/wd0ePZCOOA4KCqyWqcxHvGYwwbqFgiGx9qbSyAx+IFW/fcZD0S/+oEty5P5XotPUfwgPuF
50vzO4LChDjylzuaMkld5Dbrcfr5WXNpBgh3nDMSW0knOTB1TeZV3Abz5WJovawru58V/tyO40ys
BXLe2hJl8BpB+ca9p/Y13jcI1fcGlFYsjb+Zuqjm+Vj3qrp75yJ/KQRbWgH9y3wJMzyXS3Lv6d9q
1JIiGK5If1fssQuMWVPY94mlH6bvnTM/Ka6EVUfSYvHR+uHF+fKLb/98+f07SItItwJPN5tuBW4l
vYK+tR0scKvhUAO2rD/fEaPKZ9Hkd37oBzXLdxTaIx9CTBDcU9rylL5U/M74yDFETFZb2C48e6r3
LgIG9QLuMeHsXxzeeH2vFvwG+O2Bei0ukSl/HazLXHiQmlj8Cdnt2kRa1IqY3oFyb1MoG/W3Ku2w
9jC+V8JGDfG2iK/KPWefTRDasTjAnwbSa0ziElJn9jBxjgL85+foDCtgkXo+4ImgyGrIE+cIloLy
fsqncCZDSvKXdLgAxWB+R6QdC0Y2LIC1unB3/BVKisboLJKWVu1Ep0jDP36F/AgG6nPB0Tb9lM+E
akvszTKM3/Tyz+CdLhLk0SFW/OmxvrhBljl1dG344KPYEWBSbvHiOnUYUmsw2anSJqv2rdhBVfuP
UaFqljJajWXmPYBfFepNsb0wPw6VK6iXl9XTDTOofywW5wnOj3d7BpeN4IB1pPdExDU4uPvOXHpJ
09gFDD3dupcSROaeUee/LvVnugcyvIYLqBuwztd2grcs6YdDULYfSusCvS8F/JftrnyzOBS+lQwL
jfXStS4Y+7ByIGuXLOWXAE7RlfKBqYj7EP7o5nPm0hMbcuCLHPP/qFGyaNq/Qv+7GRmlIQhzT2+o
JqNiujtBxMRU/jZ+dIL9Gju0PECzYepwV4RMbCaGHd8AhJn34kFbF1ahDMUaHH+sd1rJUp6186z1
cfn3l7vNXaQhibeq6wkYKpJhCDNPaig4Hj/Ew9vcJuWIIRIgGgOw+s/VRo1A5xlit3M7Pj3lEPfE
wvVvL2o0fCxFFp+2j/U99alomU1YBLNWL33M97F4rRnmi5ge4NLEo0lENm0jz4Zz9x4Ot+KbB3y+
K+Ye5JJixJ41VgvI7WpUQJ4GV54dp7rnr4aDYXM40uZX0iqAGuSSbxSR3/FF2q58ItgExcholjPc
6XixPk1ffGnRxTEZaoc0Xqe6AT2n82so9m4dKvGz4RmHwXZM2qmLJXBh/xYoB48/coRJjhJRZ3NR
k4CMJyjMBhp8dReqTR6PLHbTRzensEyDpKQ/QPdZwcvbUhFCGkL6Id69kqDk7zU53DOdlJpyCtgi
2kmXY7GBOXhZ/CtcuUBMpXRsBKvDWNTLsWxTnWtWncb43BcF9KT7woWlCsXTMlBkD0k0a82FjWao
YV5Zz++x6tAomhhCOwdmv41hRQcdQxvQGf21LDCrVWSpI+XsbljYv3SUoP64N1SfN7Q/gDByvHWD
vlZIR1yFyKEQZsNdIwLkcCHyenDxh0QZrZFpEZJJ2saBzq7RxhzIK4ojdEA/J73Nv+pO+rRUOLzX
ZHv7ontN8tp5jmiDPfeRctq1iEULfzyX5mQM7CiwyPo2l/Ox3re18GVoK48tfrY1SvKQN8Z5xt0a
da/VTS1jWKCt045gpHFKylvOjj3jZLWXxUtO8R+D2LafaWE/VanW6ZeiyG/Y7+jFJ3xaRQGmR4zz
V87jXTYjYc6Sf/uWQ20DfGu5hCkKlA8tNVEGZOWvb6cnTj7z9lgZjtN1Bsxgrdnjiv5UrQ2LxAy3
fj8a1KrnDGtQMsXt7o+6COv0+0emQWwyaJ0c8F5N1qCcDOf26l17xDUm76x7iWNT0G5A7Ws4qOBv
i2vJofUCwmmu0O9bAjxtpD59WzDlFs9PWkSxLsY/6g/LCwart1/R43Y25++yqPw/PHG5UWnb4Aw5
SChyPHL3Jdmp9ZPCUMFm+ET8+BvFfhKV+cwg7gACEEIbmE4nX+o4FlAHjXO7qVVpg6WjZ8wIXdIw
rFMEYx3Th3VD1M7w+QmpT+tnkXSOhscfioRF31ZN6LuHt6rViItxNDgDhLC/nvwOhlNVNI8E/FOJ
1PtF0d1sUtGhoHp2oc0b48aWvESIe00ITH0+NZhZ7GGA6fumYNXIpRvQULh52k/iQg3DYHlvcEZr
z0hucL+khfRB5m5vFWV8EI1894cJu04L8Xxgv2hVHFJXEUQlMM64y84bCu6PfpxIkYN3H0Ar+v9v
xMRlMokMyIGykie+TpUdCDOaaPX4oXgiFleI8bn0EpQH9p//h2oesn3w2JA+WYrlEu/DzoD6dM26
ww7apVYCNoXy0jiY2txydb2l684G7VJV4uT1LobCnJZ1CuOfgn8Y3UwVkST2mpKH993OPpyymATq
BfKBoopBW1vv/k4r2uO4B7i+28CLb9+ZkDItlsz1urThyZcyjfPY18qeS5QkjfBn9vubP71AIXwW
jNDa4neCIJYNRJ3Hl5WY2eSoQzlk9uhPK/QvG2F67umhinQLsOFFzmWByRvXle/KPDfq8CQ9Vfnm
c0ajzqXWvqngMEmd1leDreW1XphYqWdIAzUsevkXU0zvr247o5WapCxh+Ugv1cntTLJWDwdCL0aW
qjKoqD+qj9+Qwi8XKyEkn5AmjXEObCyggw1aeM/3rhEFq5jJ/r/WUiRcgM/pdkfdk73dl+or2myM
NYKOkxaBoRGhmnHyyP5nE2K6Hw683kncel7V2ZGLlkR3gE0xz97pLfXNv+FUuMrEJtyonDiV+5tm
tRkAvd1ol8ih/UZKxZpe2uPd9NguPj2X011PvSj6+AN6PrjWpubP+WkfdP0QwUFmbgvRrKIsOQaD
ya42h80o513Gr5fvs+oBAKvdKM6TYQrwdmV5T9ibJZG4EFwEJMNtE+OPqmEAu5EQ6VyL8eBRZCH5
7e37w7RNpPyBl3pcaqbEvvoBc31//9MVP/amowDjgqIodJezaub68AQmMoxUCJmBpEo4WTOvYzlp
2jF6QwRMHzXIud+UqG/5cca1EEsGDAq5ucukOMy4iW/RAsS8E50KGv+9/Y16Fe3TvKkXFcmRmt4p
WyfnhGemBr05Eqj2SlnpuMSWd9YQ0iR4a4a2y3XDZlPlbZjQy+/evjZ2+GahpJ0wCK/PdJeoW4nK
ifRDwcS7LDYGlW9kBOqi6qEmg9SAubZUuJFwJw6V/NCyl6n24234K75eTj2rFBv8Lj8eHz6WfYNx
HLvUl6/PDzLif6etKnTtW93+twcoexSwFG04IpG8dhn1KQKmTUz/FJn7Ok059IMGJWIn3Vc/bGf8
2Vr+rdnzji2CPUw5pW/eeg5SA31IaEt0OiJm2QDiXgpk1OKMcDq8IDtltbX/3316rub7UzfJK26K
lgza1S/9BvGPNDO6LucYKDGcVOOw36QbTLCkAQgGMrZQcNXkN8B6eArblSozWKAVI7YnOI3DQFqb
DEkzOgkpoqhcIbWjDTTSY9Yf8AXdC34iCbwb6MwXnY7hExUgiZJEuNrBgjIEUm1Y+Y6Sv16jsC5G
lq7JdvCLfV3s3ga5bQPH1eHAETc2TKiOUsSS9q8UVPR6B+GJeAhE0ArV1nr89f4syTqHKL4oo5ss
Hf4lS/QZKVn3MKEc0A7k98RbIG+ygQyDlKNZEN+HWaEza+C679/rOJP2c0X+qw7EMbpefAgEKhuk
6QEzgKH3LFCjWpAcJLJZ20xFr/FF5R8Dqg+8314uNMi5gzUP6vrG44yIXIoHzpa9/HJ/a1Bc/a3K
BTfojFPO3gN+KbUg8gL3lf55zU4r7Ztqh1p/G6jIDnRHr2pT7jlSHm8YQ9OQDp3nQrOu0kq8sdmq
PwificSsdzWWfFYGO5EwHYaKLAiUUu16kLKYjBOvM1mJK20AEOT34dwEjueDVzCXrv+1rJjng1Z3
1wMR3IK4mivyPL+xS1WeCKO2m37Fmpve6HpW95MaOeghA2a9vkIJsjs0df6R/LrUNrmoeFrLj7Kf
Kw9Z4bKaUcf1UhFbJfz29H4I4+V5sJil/ItUbyg4ur8p62pS8iNcTvfMBgxGkDVx+L6Nn1+zNFhk
xVpirGoFYnUgd3xlRQqhmCAZjWbTyopEAqVY8fCMNuEk2JCz03o9HrWQYFVYEt1iZrm1kJ+iCKnB
PlfF9Q6xS8E+8PYGHOGyMDUwrMcOigPau1TIYt31QrIvCBWvn4CSk4LDTYOS3mG6l3jSXB+hH4pb
tCSrB/70a9S9VKsKrCJta+LH3I+1M5TSdjqBP9Q7NtGfOc5+79+G4i6fPorhxr3oHMNr24dVPjdk
TPpievifcvKbTEaNwOG9zJghCTxB5VNmQnXy3Z4HxbBZtC1JRbqh2VIaDEo8caREjpFmYLkQQ6pJ
ZVtuLMqHQujeFEJ6rsJ35yKEE2bcYP8g8StgBKhfIn4Nxk4QOIRmvKXspBAl78g1q9r5RXqG4b7N
vvECWzHTboKqIanVae/wo2iCdKREsn7TjctYU2Y+K9ks0xT5qzXLjo78qSynAPZAzp/NZYDfyV9g
oVmHg6E3RXV8YoiNLNElS4dQIR7fpI/p5oPB5Qkp7OI8ORI61dG70GHWuB5KhGng0GTx60iUZmbJ
0bRyTXDEZFv/+OIDd6h9TiF/tvkTFN+K3KrGdQBgvg6hzwUEZ8qWdPUi0jkTiWhjB1ZSh8ylD/Pk
0UYdo8dFnn/xcmo3Ai8VgWapt5gMz0tj6saN+axR6DApaWNX0vEDg2mfs2ajLU38UmoR5FRC0acv
Zg3Xgw5dvAZOigAmg5J2EbQe3u7LtmPStDP5Ak7ZDfmZNUM9zqXZKft2WVnyw9uPCx+bTs0jBpgM
eoaJw6yhRFilLwCgxDGxdWin8O2wkN8/SCG38ACWbfeG6ZqqEIsZtoc6ZD6XuukvxF8p2MXHG3Na
3k1nqSkUqpGSdtx7Fsvh2E1RBiTHjxrE4rYZsZu/pgVQJeE8aQiV9QGXNIsrMHYWFnK+uDQ+fFcK
JMn1oZ4dCStaglPRVRIFBlqZwmO+nqHoU04lIF3mAAHrngOWaLtfvvNJvUp7GEeo1tl5Q6dExWBe
rEipfFQxDmNRa8/Z2X7L1tlQB5V4D91rYvqIq1dR7ANlD5Fy58vNpof3bgSVBCjanNb7DoQC0dS7
KObIF1U4MtP3gIs5tIN1x8imgh5QYraSQ2QSF02Hc+PfGSzdkZdlcJSC3jLHmcCm67u6rJTjM4Nl
KjwQX7TFd4JoCIVMMygQSXqDPbtUnenmmGU6AmzJEz7ou4T5ULy3WPb7ZGH0hQsDo2OhO8D/+mOu
+bTuziDkcK2XO3XlLQ9eUnLSoAruvYEoxGRw5Xl3G/P7vmUvklNCSHW5HSsEhT6rUpI7x2PJfwU0
oaz7ryLg7QZKo1hUv0DkGUobwPqQFnOgi+PdV2Df7eqsbtQosNaeGV3vkJmWCG9D85wZP9YIVqEf
OU72fezNQMsXZAoLms+Oy/H4Ns+juA3/h/YzClK0PiiQG7yoZR7tMlIrvy0dEXHTD241cQf0Zf+1
VuXE2YJbAt/HQQCqc3jbW1Oq4/ybXAu77sxNRpjA9CWzSCcHl2Z5VXuJkbIGqYfz1KE+ZbRFiwat
XTNYaroEs87mG/QPkPvE2eSQAX2fqZz6+GjDlue8aOF8/Bha2RAX+5ftF9/wpnmpVzLAKthhK5gF
jPCNK8OaiOG+yXizVK+jk53z6wsHprXNoSKlZGywEfw0QazImOZx3Epsip0Y9CKL4A9aj3oShqIT
rBqkZHzCdycfqOg+s3mHjbXaxgCtUO513KFGGb1alovZheTwDnB3GzyLJ3YsNWEOpmysM4f1n1Co
YYetVTWVNTli9znQjxR2wGoy3++YE2Hy5nbk52szkug70pnX4SD1FzqV5owawztJvcfEGLDHqjfW
NsYqud5AluIEIwa7TKpWCf8T7H7farn86oGnow6LJmkdCkF2gqXmuxsA4ZPYLBtIYWNZKSmLUz89
BZchhjnnNlYYAol/baw8V2gr1AieT0bdQDHIs+iBVRQat+EbD7SJRwU4yJvFYjtH55ZTtnV1UmAf
ll9q7ahJx3k5IMh1MQu/2XB89oD8EbAWiO0vLGpk604XmD71pbZWqn/Dn2ipnea4UP3saC5l5fM1
mmj2WCTFHAIZSewWbeyyEZ8y0aDs49ThFRPBasJXjd1g1V3GCGVSoVcNckJwhND5O012U5TDAGXy
+JQsH+hayQxKeQJZ5TKaARtxgbqIcxpSYyZJZGBDSGjxWOkqMk917rV3Lh7JmDSjH/By8AozRAEA
/ZoywaFkEjMvKB4iRFCAcDkFER0ZTeFIMITqajII7yAnw3LI+YVEdlWofIxPXtgXMwul0vVSH7ra
eOVe51z2PyinMj0oZ9JKDDtIGvJ1wB9tcybKOpPTtrzoXHUffZr8REwRpa7tusBbxNicnaHA5Lwf
NVPw6NPQlGbkx8CCoK3lQc2enKs2IPUBwa46GhYbWMTBr1UXzfhSl5swe3Ik4M+llX7iaCJB3UlG
ELYIAsP9BtF2BjKNSyhpAf/9kiX/DOPEFkAQpp4kYQ1lbdvY9tvyBt928AybUjSCwNhQgrXJCrZB
kQRcZQN1sdIVVWXqLuqdlS+KNOVvranhs/eag5gJuceCC4NYCRjNdAkzltP5+ffnSE8G7uTkWFK+
g0VUsUb+m3Ns7hzgX/VPYvzL8CW4ELGUnJq84mSy3+O3gdnxe8lLt3HqzKwJryBoWcw70EUUCOuJ
SnsSr8F8k6uFjPHUtSlv2JNDpq7BhQ5ZFFDTPpwGar4eHS2JP98S0WS47goZpDiokxQqT4+s6tKV
t0hThzZlrgNY4U5H2HKgi5BBk/Ci+o0Tw2xqFggw6KvqrqX3US1hdhLKQ46/u2U0I4P4d1HW6Fje
5D+7jJa51zoNqweltIzfmx1ulj8oYdY9ElhG9I/wfKrWUju4+Ivz8KzZ/ZvA5nbaPkHWbqdkUnZy
p3rZQ4rZgjNsECf0HBdCShed1/GmZckkEeKZOwUXkiewcmwQwifOrbte/adlQDdlXlMtx/IKGjjZ
znNQUe+0SZRG2c2z9vMwTMs1fe6DtEasde82QFqPF8yTRJr1rhcpbTOOLP8gSQxXePbl3a8T4Ts3
Ora4jBaQ7jCNQMHqRVNuealwwa2GE4OkvU9rNY2x65W4Iz91EcqqrawVsfJUwpATrgZyCcEN0D5b
xwFaxYbHaO5ec4cAedmjt4nIlzZ/wK+JMRmvmOMtUijYazNXaRjgmMh3r+vbLQJJgVLG5G9fdSvK
yi3+A5z5NrqLFcJrb7ISHYje3KF24ZdLOKh9MTF3OdKwAcmB3VWeBl39pvWReyfD79TtSsPId5hg
UdKHvdToewylIlJ+RaSogqsxHwVwT7xuFd3XLG4A3Tr9lm/nwmpwgKZ90lWFW3EOfGxWB4hKniy0
pqLPDY81/kS4Vh1sLYwF+qRH9sQ59tliglWvFddv4TxGQAHni+8Trov/n7g+80wwMMZRNQZq/bVF
5dgGsacZskOQQHN65L9WdNVaZkIxSPznBXlwk6nHMFvZjdnrrnTuuSx/jxtElvI8RCqNO1EisEqN
ZgpaSQolBIp+IgPQjV2GoyB+eKIJKiaYuMakgDmg14VPEbyHVwKxs5XeXJZm1UiJFl7mbDCFlhhI
yGwvUzYb0EjmJEaakgjNC9Z5DorN569vMU0e39OLuhtu/vHsNJE8oFTuBsXMmVZhUiMwAnjRtC1u
hvKndcmosm0wc0qFesJ7FPbLnsze6IHlWHCdoZOR6HlNTaFBBh1PiqcKdMROntVRoZ6kyIFEkxRP
eaP+8IWp9BctUHqWQd+uhTJrgJOSBk2m0xA+V3yjBCJ+DDKukSHjR4vtVxlgrco6Yo1lyPvJZ9Bz
tFmMuK8/5tdsIws5GSwyWPhRTbJ59sDNWnM+bIfa6oCfbGm+kFnVPjSVEsuN4Y1K33+4HAnVVGx5
FcoaBH3b3Dk/X8J1ILqqHK+LR+PLi7Y/Fl8yS5kXfw1QR+Kq/xvXrakAp0TeYeyIqnjaifSaYEXR
IngtwaR+dL8M5W4pfhE04eXH69n39+XuFD1uwzgzc2i7r0QIoRcZoLAFJ47s/CXkjUaZtSLUXEn9
pN+RmXpSC1InXliOhZkS1bUsGmAj3ksz1b+M7rI64yjzVQn+jwtauOc2ahXIrCWbpa07RGzGyvzH
ATHlDC8A27Z3SrlpGCd3yMDBCPWYzxsA6kc+FAf6/IzyPCslT5G3YshQkAMllqf/vP9AtpIaqMFw
NE0HZmc1d0zuwi7KNvpeCit67YJjhwkXdLPSygdw0WT8P+/1hXu//KiYXtsE5dJZ/lcpU6h5sxP1
Ts+/YValJk3d0NrfhtxbFwQiRhi48AaIXPzpAJUVKjj8Br+Os9pr6H7ArvoKoAiiEizB6fQ0PTdV
vAlpA3nyZEKWZubTpHLKY2RnHPPTji4QPQknXKYHvBhWORSh9ZlttNaIubM48U8eqh0wKiiHPAAI
t+YPsHyp02VvA+QyLnWbSy+MAXkLO92yoxpIN5Nv9NaNBBl/8T2XWiLgV4oW4ALdmuMGNBJ+it/h
b5MzK6Gsin+d4RGlju3lfpBMZSTPKzASIq4TQTGyPcH3aSTxvX4qVHx3ez5p1e/48AKKmSBmb+Qv
O0he0I0Jsu4PHKJrqO6x81HYnGlWf3PuTGZoEC3pYCOy34AsiFaXp9Y585yRBSdND53xpLBeMKQS
b0wxxoDwa6X+FJxTwogG1WBRRcx6eqzaBvtTE8JPkS9hGz0ZPmNSCBxkXK8DaFQdUONwHwf1UWcv
5Couxo6fcPln1nVfo5loDU5bE2E4mqYFbxrnJOke7ma9w611Mop0HYESabO3MdPOP7tr+fJg6cgA
Amrap4XPHpMDbcmIjkQ6enW3e7e5mqLdLp4v11q5uXh9pUGLN7IUJyALU6XPyOeAk3Q7x0zx7XLS
P6r4/zSUQ2CXTD/7oKO5/yEnZOBwW2SDO1x9rH81HOBK/ITNv7m53H1DON/Y4QfyUJn7AhRO3VuW
iXDUpq3O39mbrwUPY13V0LWzgHI+xrbco7CQYuWfnUYQhgtpSO58GmGa67KW0cbPh8Layh4uAf3m
PBmzXACKloK49oDOq5K8TOZpIQ16pNYXDum6iybf2wW/wVUaZZRujJei7UvrBjtHqxxohGSAc+Ic
DW9R80l5Z7ykKQOVO4lDF9CcQ5G0q3XlFDcJnIvzUqoD/JbOP6TS1Y/Ugg0lEleWklkOOVejhmAR
g0FlwY9NvjyoBUTErueDSDCSF26DKmLqPcSRF1C/n1QHZ6+QXswJ3+lykUetwUJFD3+VGVgaP2wr
kqg3DrmQyv1avK0JwmaXmZgEib1B2aFAO4zFP7ABEeYHAsUfJfngUyd+6wqM8wEd7cssQiyoK+IS
ZLZ/mrVsBdtopl/zHT6v0BDQctxX/k58Yhb4vkCUfudlmfkCp1nR/N/POXEK/SkPWRnTp2hs8dK8
IenNkNhQwFCXgWek+6p+JzRJ1fz0uztX/4TuD2lxFn+4FP25TdZ47Fc+dK7c8tphwxI/MuZNL8hg
3qDH0BtdgF8MoVWpT3fYTqriO79F4t6maw23yFQJMpK0uHE5L2hg/lCrSAbWXnTjW4N5ZDe2AJj3
TX2UMIRO30FYBai3sCe8gqifsnSD3JfPrvBpB/kM9YirO1e7MVNmK7sP9cDAxcrSYu0GOVzUFn11
Othr+liBIEe8zuNo3DpHLMphIDMyAUWVMESo5vJNYTDiA7ajeiubb26pAyrQp8XYKAJuhutqghiq
ViUGEVqXPhoGoZqEQEKDP132dwcgoo2NtGJCyuRiPoAGWZYCN2wzhtWqd+Q6H1TOVIOZjPnvNX7Z
L3/I9fA1vI+yD0xipcebVaKGBWiHMzgfoHbeB+Ro3yGRO9EuYYe8Xcch21uwKBjBOAwhRJKnlMvJ
pcnG1D6v2rn8hFgpbOi44vzgjdzkMDENqtbCaRGURutPDjj7jkrUsCEFSrYOnBA8FJagNS6GgbMb
cDkdeXVmlTZBTFyDGJO4NTjkgGwQ889SxJGquRPoK1zDDQx88AuOs2AR6/kootIBAQJdkO08q+Xx
OXptImszVJloq75qHlgRXttpgKuuSJXOObq/XoFVxJBBLe8OlmjGrOz/NsVp+VKVirkXcqjWMcH4
8fnyU49a1WFuVAJu1Rkb7Kds7NP5dX2kwz6eFgFkspV3JZmBF891Q9tYLK3r1bFcJxwHCjxhAqeC
3Xq6+8u2MvUTb1GZkc3A2H0g9Jk4b2XgfpDiLEVkcW4e037YYqughT5IvgBsKUzbhDbfUmQBKRxL
rfIDVuXtLAia+k2aJdfTUeizkVwnO44z+es/M+ONmlAiLsSnaf6k4aaGVDGY5OrZn0VOkjdwmdAd
povJqJsO9I7T2vrqA0t5rpNCaQQfIa5RDDWHPNztokmep7wS5drFMDMGcflbxgd6vVI+jc3RSBoX
xc8VX62EoYiqrEXUiFrT05z6lO1fIq0xNve1KXOz+LaEpnQfbmjeDyTuBXwrf4oTd2nYn3R8w3wg
U9g3din+4ejhxWfLwVqoYU2q9PQmEB6IVsuyzHt5WB2LkqRzsvdLQ5aBiaHshJzT7FTIgn59Af/M
XJayQkqcivlTBSBDIY0Mwu0HrJro04YaxECzzmeisjpZ1+gVngN/UBbEyX7Lqfsfdz/NjHTzpERN
TmmfQRypaNH9pAI41rdYHKuyyjygkT2PsQL/j0Nk2Db6rB5MDFY+ixkQWpL6jCEZ1HYotsWVyS1u
gKa7uiKgFQR2L/rB2AURPO1g//drsjIm4Uo1PU9WHyMmysJr3qos38Cxagbk7cYnpvIX9tbHDgWr
w67tJH24QO49E0thZsIzOE9hjvAY7mPa5BH1VLco/srxV0xd5vV0pppdAh6qafdyiQNpDUKicQ9G
ee3uA54M8KHiaZ30sR85rVUr4faDeCW3z+OcxZtjabpKlfQYRlUneHnbKdFvg/+w1cB+anjehnR8
eqbYq+BNfURW8rRqD+bVGFelFW4mBx1SZdThFCa3szIfoJmg5JDzvtl+9MvI0Q+WkO51KXoOmmmY
DGz6q8dSGqpccOPKOpeFQ5jhpJCES5ERPad2XqY+5AXlNpVo3WYRegofZPgfIy/+/BFvck3Czlf6
7oK8NR+a/bS9mfjn6P4t36znq9KdKFtMidDXds/lEx+HCT0cOgeyzJnJgNBUj4TKj9u0BfJLi8ra
oGKrbowMV4ktL4K6PVpdaknjVTbIF562T3vVRcHRqxtOZ2+TfAMwd03wmzTC5St/K3zVJdZ8+n4f
bkb4rY0dgy6IlzCYHsGYfDwV/fuwC2BoRYkSJbjBTa2aTaq1SPVWhT6PgeaXRVFNSgWJwFQWbDme
2DpMD4iY0/9C2/ShA11PiSENJLf9aCs2v5hgRnPox9VcbidU+yU/8fj3j/d7d/vWpvwUaawujhLZ
UuXn8BUJtYYy0WYmnCRmlNcixWME6VOKpKBNUfGP1DmNn+dpBAlrLGEkT03GnkpntgjUZsYuN1vP
zYktZxm/TePFyI1vka+iJ0CbrFe9uaeGmSGyqch3Fhu/dFkg7G01bBq0Ivf+3kblBeq1narwQ78+
BRiSJjy/XrG376bP5+AqjLydEmxWriVejBk/k0Pe53E1zguxff/+pNalth24quP3fczJK484SHHN
WM1X4pQ9ClWqg4KhDA5aVmm4i5x9TAYNyUKenwNhLbbef+6vZmxY9rfN67qk5+DGHh89y/v4Ftf/
+7+A8aXfhjoCnQcqnvvaUClW4nb6YDr68WUeruz5jOaC6ffW06EEGy+TgtxTPeSgOgt9ShusDRgj
KUODmXmh0Y6JyelUfVttzi6wB+wL827XAI1pOtZ3YNIdj+/1RWeOjgDEP43e3NT31zfO+4nnVqor
uKuqyE33y0HzSJjTPlrJPWaZ/3zHYmMjoI8Lv3lhdXVJwkAAokvYggg8KjPnYwsjOpeWCk/Sbt9x
tVNwaLKi1ZZJXd3Vpc005MMtW9ba5q4D/dyDkFmFlBG91mDAU7GzM4473SeEbqyj38ho/CQ/k/qb
c1UqHXIM9j0zinU9QmzFe1Cw5FNeo/54BKWSSF3MTSaR/x9mvKpA6KkxaYsDv08v1B2ji8bz0+mc
MkszUdL4SksetHf68T56etrYvt9lxhF4PlcF5BzM9JQ1SVM0jVxW5m+n3Yk1uJ0paW+WGWUG5PfY
Z/CJ+Tpk+fDwBLEEUheq9b8aj5ypvEEJt0mrL858b/kvf/Eh39b4Ak443lBadEgP0PclIFaU6nK7
UHtCHoSER/oTgy+KMGXoRr83JQaKUtmh1xqSiehtykTOR/BcyzYAefuB/cTy7DaTzN8Vb4ss0pqO
aQErReeobzsHnQrE8BeWcZV70wh6A6w+Jhau0kXUDVZ3P6EZn2tKHXWz7Yr2G9eFRBxc9XqBwRXc
yD3zeHfu1ahO/aaNZAwze4QmAr2QhWiQqrsb76B9vrw5dGKmHHnYJslFzEQ2oJFE0WU726PD7E0l
Am/Jn+WOjrwCx4UGKw4N+MngkDZ1Im0rJcngWvbEvQ15fX3p/hfvo5occIEOCTSU6OR+T6lAZecP
I6reMMRJhlO8H+kbb1u6k3wXaC0FGlXQrmmBBX3rWBDHLo9rf64cHxaaYG+hWIFHEiC+Bnh2P4eS
FSFNiNqCHxXcuajs4xBZQh3bWdf0FBw/QBfpYpouDxbWrjbiUOpK94flT/aSHFrrhInZgz0pgB03
1vseRAQX1pwzBkHdctR6Q+ho8CFQaWvtvATunYXrtdvlKsum53AMRMz7gdLsxEePHMKS0nqVjdRU
jhfkknChB0X80eiOimyHlS4WNyqFioxjzcbv4MAKeVeBt2M5Nritl8Qr7vS/0pznGDHfc2DnzFCu
vQ56l+gfcWJPOby0QD1+VDT6TLPMJ430CXjOuFs04TVql69t+m7nkePU+zp9yPHmJ6cIzadyx8kx
piSBaePqcWh/ov8TUAVKvAunHE+Sn/HiCGbsRb0Hq9FynL5mA1nvCwuwhSX/Sd9JDaCICM4nUJgx
ezEeWgRNTCbIfl7iTYpanFBxnGuMSbzbyBFb5NOujtykk4BiyKD3lk4ATSttSYMffWM1gK9zvQ6g
by8TKNzh/vC89UhR3ZFLXspsdiPGvnMFJT9eUDgtxYFA6/xcLys+wOr9jL1U9NeYRwLhbh3QGQ5i
bjgFPJzlce2e9c5jW5IiAbmz9crUy4GWseBGWf5YuyAL5SYv0m1JABbrEE+tXDPZrVU3WTpWTvEG
m3OXo51U+fysmyhpxJRDGKlJb8o3Rf7HIDkd6Ep8W+m3DFZHmKI7Hzl61aMuz2/IG/rX8eglE/Qi
arg4J2xmpAbnwXAgnKJBZ9s2tZbymxLDKOJXKSMs1OZFL41/VBhNV9Z///nPGT5fVcZRg96DeKJe
2MBoyLAoE5oHymm8ODc3flVKC5hUcwCRppu+x0Uus9+cf+zp8PT2AsXpWEre8TvdkT3aBF9wEXY7
D9T/eobQU+lze3wvlgjUApraPyrH1z2Bu5RT37yCcEu1e7qJi0kcmGoJeeGg2LwbKTtTBOxW7V/b
MWhHifYWo2I+rX9dYaeC/0JvBWyjbggNxseU4pS/inCvcmHwdftn1HQ7SiYqMeALs0FhQdpx2pth
lcPmNsd5s5gGkCSw5agry+8sOwpqILCxC+nh/o2BALfxfC7cI6uqseQAx1WFSTWgwhposmbvQJxD
I616VYjU6zc6jzOxkzRaiLv/ZBOga6rSM+tgIh6WtIS2Met/yG3tgKhSWGmNwVrnAhevkHDNRKZq
2IXmUBT0QTLO/VAh91FQuIrO51liWEdXc0bItrgU2XBOnJe2EwwfXS0Y5YK1ESaWw8YK1w0SEqqZ
WGV+YcojOzjRWd/wXIqNGPPNoQOz61uDdaJpVueAvtUU51vjBlEUrceQk2Ow+wKGMANXllH+GTXn
XkFdMBxeZjoRmliyHLJmXdmdwuXe1OKTO01DU1joOwnxvRGyY5JsJ3RyliH5EmmbMe+D4M4V9i7k
LQ56lhAZn0iDnEvWxCEW5E0YwxTBPGZE+3pvhoI9q38n57B2LzqE27U6uTzjr5UxWj9H25NQYgXW
kl7j8zcQ/7gnaKBPw9PPvcB+JHoRmNdDqmFqOXHdUi65qkd7LicT3ohQmyovrXgLUwSoHQhMc4O6
MxvkCLkslLVEwmaCIM+izhSurWuIE6sqh5ijwHq+kuiYnNl5RB8OEf9xF6h2HtgYPu8iYV/Izcmn
YwdzjK0+19KSJkHv4OY911i3Z1V9pOc7fYxNRMqpcYeDlXI9/eAoN/Ewg38STHvnmrAr+DJgKMcq
+KbVk6+GQcAB4O0uo+Hyr8A1oduKMT0Xx47nOMRHXs5Wwmz0j1pRCzK96kbiEFtUaT0l6nLbnRkM
ScrhulVR1E8io3HSSftch1nns10huGIc4lccDuscMuMAMqMPgI7CIfeuSXVvUUg1Sz2wEePWdpFS
87QJr4e61jBP8kkGpVVNTdTHIAi6Ci3LvUoJibXjmWyEU5WNaZ2oK1S44/V1G+uwOkGfSt0Fauro
M7fqCGW/3W9HxHc6vTVQy2vkPRbrrqETjvF4MvlmrfEJ0jQqoRfpC2wKG0YeUneF+uD0QSThUPac
rXhsBzzsWJAAnv1jE+HqRXEjvS/vTnLvVPsLoXzMw1t68zPSOBXxwDhsCcpw/B1hrqnGTiUNwtHK
po+VMFl8R7qIuxqOvuBjJDOVnr/GirzV4rv8DsOGE98H6UkkBwYSreXNM9qd9PwDl6jdgnjhj3V7
C4shBui8mLg21oX1+0qVgWZx+G/yqCgJ/7B0sdQVfeUjes1Ljm+fsx4q73WRD7VdpYF1IwAA5VoC
+RwtVXg04sSptKMzAuz5UtFsdvGgoRrAIXxFKpQL/Rls856QKn7EgWGx4HJKXOjwr9LSCvsovW+q
Sl3uMG/oPPQ8s4xrpNUHLxN5fCT2i/jFl1LfM84WIM0SyTwmSPhLNWqLVNndhyiZhUbwqH9VjQdl
Tky8E1bsuKDiEYsbThs73Y4aXrdzkMqmdkI4sCQewZ6dMhrYEDksUxOPU9748m2t+pf7j7/l8heK
N0qGFwj0/G7uDkGMUyuw6CA9qV0eyUODF/se8681hJu0gt2XLkvUbwd6KCiM+TQMXpAM9gXUGzPH
uCxfmoWIZkJzwYfBhK4Z3OYmg1ElnAkNwBhxeyPslENWBLc+XP9MHEzGQGa9JdK8l23nRGZcyrL6
Dy18BvwAxuiQpAuJWyZ4xZckNslstJMNoad+KwRYnjdWKZy6UaxBzq13Pb4imSMlMdlTmijuzgfl
XJmup7AqZxQf9aeVbsfi05DQDl4tO5k2ghWgVThHF7qFDXAM93aYS5jDVeyGnNWU+cyImocyDdpo
PKWf+MhZXQjMnzrxqTgCKtikb+tHV7q8lxj0cOCZFMPefcvwXw5urrLGQLeO24ASBlO/oV44TPkz
EuAXOs4ISClI1ahRi0S/fBT+QjuLKeIgRgsjAKIfFb4ywab3KqqYd3ChwN4NZWNbE6mwEwD6SHPB
0il1si57/YJdKkm6rn2IYJTcQ/BP7qFkudjVOfFk/058V/tDsMXph0UL+Y4J3+Uuirg+EgD6uYNM
FuFSu7o2aPeYCTGXC2R9NzXa+JHm+mG6GXex16Az3VkXpTlI6m03MlHiN49BWjuaSl+VodliEjm1
4x7jPrvBUpXZWG+FoQRLluWPW3NI49KVWv3YEcSFDitVXjIY9FAFgw8zWEp3Zj1kWTnfcfyC4KS5
q2Cq59FdMOCPjUwLMV8x1rw1kGujQbVWnX4+5KZZu7Of6dX0R0Ew0nmFEKPABRw7/2nKmAltL4aj
NfdQNKFRhA7oy+l1p0owbEmn1qccZp05hR6M+fIe5ilFSeEuK5effu65d+YoXJrAAPN0IKn51nRt
EZaqxMPH8YWjmyOtgQIF8httYOtRUOOBnwWX/hiBEr6D+Q+T4+JecTMJs7krgyl5d359119L7b8q
QapVE10B+qUjgdHNaRbgnLWrZge95uSrh28C0d3MyOm3B7myXwBq7ZkwJP8gaHOicGtR/LHG8yzS
lFE+MlhGsPetY0p+VEIp3Q5zWsuOK0lttGCEdCKjCZPxLoe/7GdVUzl35VRHDPyLZUh3H3WhSOtz
dHmSAFHg5Acb3FL/0W7MGrdejz0G8Es7bgPsW1Uj7ZDZvgwkHo78O7eUn4m7G2YtymPMC5iU77sV
SruP7DA28Rax6Wy/1H27XhZdW+GOfZOLObuApXuB7sZYB9wtzBixt4VLuX5IgzvCb++jQUKh8X2m
4aQlMyVw9XGDX4gCRRNn4BkGpQ7k71iQqPLItlfcs9h2vq0wiLqr1zvKMp3wpgBxLyGY+N6iNIP8
QBFtqzQm0NkSxggSUlgqc15rnRc5YT+ulxL8atY16jERYLujXZu4mZa4Ia4plKYTDXwdSCY5lZqq
SgI204zrZMd0Z3MOJ9lNnuPq6lX2nYlXKKx9uFAHpP4ug5EkGDeaxxzGz1m+UgVdxZu4vHs/lxJh
PwaJUPiIAAUgdRVn56Z7FOT1zrT3vf0yOZBA7r9TIVy9azcM8Tyuz9PSF9LAARoQ6eJxq3R/T0KW
KwBwRKKdsYRPOpZPJOWDq63PS5jSgydzQgcwOb4mJOXC4LIItFdZi2+3Xu5RNUcuLQGm6hRdKHgS
s0+U5E9oXFHSbYIdtLED7Nn3vAbX7Gb1qEQmd6mLZxKOR6tM3G1eByCCny0BQ4Bqt6I0L4dh0ERx
b5mo2kVtj3LWUjqRSStGnSUEAVtpmXmjGJMCUhmiitzCjLsJGKfTrMArWgfalxkdbuN7BsDje625
BPRmZ3JGq0TPjHzXwTiFYw4VDscm0wedy6Cjwhb5W6YqYTbi+iGVTaBtZ8MZaGvafUHeVELFvzrD
trxOvbpPlHetpFEDGOutMCa3MPJwehXIl9NUyn6gPbVw3ApSHmMegOPMYpYf4zB3ziPFqXtUS+Js
xGvGmnAFUDnVPUX7kCaWU4ecVvWhR4Nyc2R2DAYT1O7IFH2N8vDh5DGGC/6sA20ClHw8Lmr5wknq
nEVZHMiPU/wT0b/d272hylUBgRyMV+WmStyc4m1HTo++JU5M7ADSbQIxG/kH2wELI6nEIQM19VzF
Yj9ihvIm7QqZKg2sSFl5hfo0C24T9WZSmzSVNHo4uhu2X1Tqyc8mkDTtdtutKMe5t6G5EGAaw3Z5
rvlFsDDTsKbfuF7dN5TO1D7Tyg9AsH4k+PLeBJB2hO/7c3gfO93F1+/zm2sj1OUmoqY6wN1SBF81
czP6V8tzldGP/WT8JvNXUf+FIGZGyfk2HQ7xDMpjanNADEfb3xNPcC+9Z7+NkwA8cIim61ZBqnhv
xq9T1vL0r7Fcx4jgW4azAqdAf+9VeexRs+eUaY79mpkatwBqFp3YgK22+S4Lx0Y/+06RuzRjJb56
7ibSrYfHXm6hGD2DWmOF/6PKQJoD+w/lahEDf9w3bAEdgufy+jASgUdj0TEJ7RUDbfb4cC67rC9J
lna8aTpfUS8BHpeDobkiKoduFX2yxMMvuhS70G0bJCJXKLOL9ycgoBUqnIdi52WW0PspcWX43otF
b6P8B4Dzz/emSPUAOJP/H+XrkHpBKWO3vEIMkWRRAbCyGmPB4Bz+BOQs+968YRafmJyZWJkZkb6R
/Ed9K/xpHYNxpAgwd6BU77UWk32JDFjDI7P1gKuECwY9BBuemIqKBTchM9x96fT5XlRem3S/C1Nx
IvizEXzW89R7qUbjfWWbgYkjJEa701wGdH1B81zLm907aYkdtSXvKWd7GrJZuwpt55BOowLLg9Kt
oreqJRjFVH0YFKadkFB7D60Ew0yReUG2GdvtK8TV2UHx6E+ZJ1hl/pDxO2v2PoXcQikvYRn8szpF
j67YEnWvTCAc9MGcpZoacE3W2ue+Xk3XAl74xcLFaJfdU2KQHgdumQuMa6sT0ZcZRd0SBBu+hwEr
qPHwCQC4sIoTBlnYdz6Lt85Lk3AqKMKY0K11Dv9460ezwcbxGtUXsET5IrYnY2ZDSyrXrSPo1Zko
ZgIFw7Ec5Vz5+7YCPCxCxzyAVjgwcWd9ZCxbhaQ0Hw9NbGm5IVUte1b98ggnTErHkrFEuqE7Vcap
zeqziqauE6wOErXThE13Jqpf4T6PAsMdWYZiARUJJD3Owybyef039/cV80KuBgyZlGLsKwK9AEUM
ieRKepTpdmn0NrbH3kb7n2NtPcp4ZF6BeNNNVPjy+7jLrOh95ihPZJOv4Wmd+4LcmAx+ojvPLsVw
YUhdAmomzkaQYrR9JTxGVK4YwUo4acWAhTJA7/hyQwIvrIaSG6jJ/Aiovj0eLBqQzuLwyssHY/Gp
Xu8IwubaeNaj4uk5iJaF73tYsZZ7OUgdrADccWOT++Qlxt+TRQSb0k8DWSBF51yLNWNw2csttKlw
+bKFpID5E/cEqZykdTPsLN2YnKDT265I4rh74e6lDSLki0ngoGtoApalObv3hzWvGEcbjUGs8LuY
LjnkzHT5dlC5ZM6GHAd8KcVXgCz+Ms9zCqjZPK6SFNYmos4xXv4SYUhca0H8dbKcbkSzzB3C4mBT
5unN8HdYOC8xU4+z64/PrueihOu4dpGXMlmhs9XkAM7CQ4cwkdaTlNuPc3AztvYxUX99bWZF5/VM
18wf9U5rNrVm39w+BOI4T2iHW9lBPnmdoQjKgs/nhwRXTdaORZQT1y3j7qJKTao8iA2Em7cAZC6j
KagDU65MvVbh2t1d6yT93YRQTmUKfAOFiR9W3Mb240s5+k9/mNYsvadaBe7PHWK2hJ/811e4bBcD
RCrOlPT0hyhZnB6H2Y3fnbqmATd+qLnzmokURkZO3ylG2miTpBlV/L9QSE5I4ugIPBcduAcBbUe2
AE0zoyncwG7OhVMpYMDoZuODhukGaMBXfnUUliK1yd4+bX0pF2FaFYAlRDiYvu2g6+HujOrs0xBb
avEkQIaVSkwNl54bmSy/MHVeXsNpQ+8xMIhjHJwqTYbdFPZz7+qFPn+XEyD/LtH4OU+xuMQAmdlS
2nPLEqH/9myAiyugWYbvdCoxXFt71AkAdvGWTu5M4is8BYkcUNgJuKxPaW6IQa35AMrG8c8UjTqy
c2RoDGKF5NMJzqBfiHZxjctUe3xRyTHZxrkTl0wQ8PcHWNOvJqSAwVVWSdMcI8E2i8TmlUGGgfNE
oP2OTRLdvdF5z3nx7nPuPxKiEO3vx0yQCDhyyR10aviJWtUchjnemiTEFPk8QaFIIlP/2u5fiRod
g2DPr1NIvrm+0gyRkr+NfwsfML8MQacVQd1a0SKXyi88191yU3MjnRGmOQOA+QND4ZZzvyzzr1GV
4oZlD8dY24bBZebWSx6yUzSZchlp2hQQzLOtfLRxqmSAUaeP61HaMMIEKXIsY8ijbfCX0YfFu0bz
5gpUP8mMTMVKCXPmGSqVUiXiQBgPUpHxbZGaRISqLdkKQAa9nokx/DQvsD3mI/CZsGSD2djUjG4f
XNTPXDSYeaR4QaaO4YdYWu1m2JH1U6u++8vdWhztf6kBUjE60Cv/qpT7/qs8kcODRlXJ2j5AIA22
Vt0JYp2adxxn0u3/YhgVtezKI/9SZ6REz6sSs2KYg1ZwHWYDAFXaQ8UUGap8W053pJAO76YN8nzx
RD5ueH2Z8BTBO40DxAEAMADYOUSj8PfEYoO3yzn5JGuUTCKJiwH+JVaaCIvZZozxozd9pbtB6Xrs
MjUSpFtVOKAnqPo4AJL/0M/kVZ4mZQPa4dNuKuI56ygSRSG0DkpNB7aCZ3cJXUcKvtdsE9ROQk2c
sSjtEyU7CwDFvX9eCivdOcnuOB2mjxoAD6SxNLaXGkldE/2mQqc/GSIbTy5zx/tQJIDHOrCx0vwd
xRN2Q14iwkNVBIpKi1dCqfFVSQwbOLr3IkIYO+XKYO+V96DDFWNJi0mRq3DQcUmkdVy9vA7D0onW
+83STEfesC51S+7m9jjSyV1zWEsyY/UnFcRH0pzK228Z9OYH1FtzWmuAYRif672ZAhfBLU32uVET
I/Yfczlrf0C46aryE14Nu2PM3sAIMw/BqhMDcwmgTPkRRvR8qfOMlmp6zP7f0adVgIHl+GxpDGDN
z0nglpOPRIeG0d1TCxGFTNsfjKbQtVxy0TxUnWgP8tAqCRvUXwWSkZSGoZUXY5PPAuKLa8ldNgCH
eSggpggB6DdZtDB1Ygmyj3CcQwdBVpVVJ2Q2tFXRgdvubOBlecoPZ1eMIzzpY/migtdgfJcxJ51P
Y63iTmo/Qw3KAwRyWZlcCZV5qIBef7La4r2nSeduEKOr1KE7KRGCtARJ8Euy60qPZf90aNioAq05
tLaRIF9KxWt8dUQuKGUhTIJr1IoVNjd/ei14JqeryAAlEwpaEl4TB3UNWmIpJhiLHBaZdlqslYsr
YfDVjS8rk3de2BImqzlhQftQzJLp141pJlZvx3YPaKfIZxwfhWkdq1KOoo4wGH0byUUrd5xWiFzy
1jN/oUcoeu3ps737Xwg/ozP8FOaBpW1992kUeo6wt5zr5/e+NKUPjAcLQJfUj4goq8z33s5+Xor9
8qXZXy3dS/T+8AwdRCfNuFs3hikb0I78xd5d39HpPBQHj9+MK+eQPRvAMPFHvV6xfO7Mn6Idmqe+
WjwSWMDsdmLgvAz0Ma6bHvs/5JRvHti4ehUamfxlFU+d6oz9Kj1KxbsVtqm+I4rigSzpDtOuiJuB
qpRfeErgqdKEMMh8yC0FFw0YTCM7WIfVNGFUKLLK0TqIOip3fAl56+xl31RTcEUmsYcFu83E4Uan
U3TqPttmhYjkxQb4lVOw0N33QYpK6q0v9j+59CKbiTg8AdUOfj/KhLmsWJ1rHh9ZgWrQ4Twobpx0
3+mJWsI5Iye/B87YANdGRzhc4rMARuusUrCoxXKL9FpLlZKIrsSxziz3OhljuQTRl/238RET5nCy
2x2oT8WeYcLkGiTB25OhgrZNS00Kj3FFBbXmp5MmFAThq/p0zr6P8yxZC85bFVZeqiVEMzwPzat6
gecD736a0kVqmkoqCcq3KMyqWShLcckhEacsQMgKaOtBbvqq7me28ZbcoO7JBbzDwLhqH/h53hNN
ksMqPzAWM6EB9FeUO6B974w9emgUU0woGNkKfIFfz3IdFGZM9HQOHiYLcNCBI6bWCKB50fu5eBEJ
KAwailqUJtwwwXkJvFojA6QtezZM15HJM994JgDy86XSnuTxlmrluNiamkqdyn1jwUkNk7SvwXBS
J4yX/F92kpv5nHUc75zdxklj8FTqe5zdtOiqmOCX+7bhNQL7uLShQec63f91f5m2ig3GcIW9lTwV
wQ8CYen4LL+Mp9HaK0fEGbHNt8tvxUgMUObPME4yiSaCJOhO3t9M3WBEBLlNUl5LYYatR8fHgTHx
/z3fKmQFIVmY8MWr1QDiEasWf7IAYPXv3vrPIoWKZ6mKe6ON2X+D+X9SXaM/mnjaUOqDNaadETWR
c7jU94APbh/C4GuKLeI7Hyml/B231PKlCwEMhHSy+mzqwoxcHEmo44fF4PL29xhwC6QI4dPDWnKU
PGa78JlzvYN1w3gJBAQYmlOPoa4RiDctYxsswkb9ErmgGio89FO9YBLpArPcEqP8Atkk1jxzlRX0
0Q9qxQ8Du2uQ0jImC2I+RiuxiZuZAbYENCBYm/WIa978za5fsqJWcnB11SixY6OqMDW6GYA1zN1p
cGYa7fcpTfApBEIS5DKaxqIyrrfM/naf91MoLSC/ns1DjYMlG9+s29oqzb3WKJ9PgB6YRGpm3s8N
cWqWnchX49+hd9HS/1IIHySi4NVZk6p+OIOmUJ6GQPBK8V3SXeFAHLhune1at5or9ZzY6Z4ihUDp
jYmIQThtBmWrfzGMckTigWfLPWd5NPZzEShLbkrqRwcxhuRAORL8NEpgDOPTdN0v5Qqh1Z6DjXGs
Z59UOV7IjW8YSCcjrgalVYkja6OgcxfkitYVuvg00QwSCiLkqJrdFOMWkbsTMIV8tKzuuw8/qtq5
gZCi9W1dElqFdwVhItBFoyvIZcQgghz8ZQGw3q8qydpL4ZicKrSLWexD8gk0MRB/SBaBVHr+FH4s
gDToAMzTjUKl1Pn2I+NNa1VAAYJzvilydtwX6cDvnliouYSCgfjLFv851iHgcf86YN25wAkSJS8z
YfNadpjwc2dofQ6g/UW1/v7F/cFx8Y3w1XlKklSGlLA9M5fyxHjLYEY/VkFlkvTWVB1FxXMg4Huv
z7ZGdqOVylrMNS27z3cknE15ozmZQwZFfSZYAAdmgkq2SgaQgr2wdnkbvViq3b1GXuaEME1APFYW
shBtyTW9MxLbGH8cjV/skExy9IaJn66vKLKHvCsc4Jdq4IumeTnKBa5+1V4IVHHpVEHLVEJcvxRu
FZI15C35DJbxiInpNIYTRvI5d556WyDxUTmFFMLMEFMNF3xnHGaCtA9MGQM2b0LzYsnrqfGhxCpS
cO05aUqtDiUEXiNDHWJT7m0SbPmEymE21r0IU6xjOX8njxC2Y/WBIhNw+e40St6MXEikj7FzuCc/
b2pLBhLQbyljDI12AFHUutDIrk8Yj5AuUuf/bqKDpugZDOOLDtCuNWMHN7+k+QMPVe7QjC2226Jj
wcyo7NG4jvWFry0gGrSBKkwE/91uEifz3uX6D+LYxdb+wPM06GhvYF15YVlnwaWD9+gXYM1OXj0x
YTz1gXuTFTaKqdjuCcrlSpBUZnIQZODpTNciOrffxUDIQrcngKKko9kG3mC8kKqg3Vwdg70uXgUd
kSlQa3llnXQD3hG4tNzwSMcqPBtOgbb60MIryzH4O9UZ3cZCIo7A98yb9VC6i5K0VJYlLpeBwOKF
by4WxkpmpKdaLl2dfM/Ny6rRtSMJyKHXNG0qgEMBx+EEHAIv/fuwLukzfF9hcXBfY1eesvY8MMil
5YbJvkyhu8khmhno8PpS/FxVXxrTkPhP2+y4FnmKQZ7b/OGWeJZwl1dMKM96ldJN7E2Xo2jXudvN
09nlHpiwS2guQIKd96vgNLgxdZKhBRa1NPURVjJRiP5edy9Or197etlv9DfUjUSEsG6AO2GEizdL
yvoRfp6PVXV1f9D40lu0pbJppw9TcCO2Dd6MnWP0/eVop9gpFupnD2V6K8Xzl/YdDnflZAPo8NWA
JkW6wDxdYK82hQckN2ZrWWEQl+fBbiPfzkHw4//nnk1b3XLqHmZetpScc4ue4ZL8FmuQbjHfXQrB
O9pHes2ou6zIbJnf335GUxVJUm2X1ajHxEA2SS4Nz2K9fEtkAqZpSukPhcFRL0+i47S+4TulPWxI
ooqcoxch+db0R3harKUaXRLfc+VIEaabBKWQg5ijTfMlvlSSN4vlz13kf5QH7u1x5QmrAoP/xnqr
2+lnN8RM3sJLaJCzhr/zvNtY3sADi2uUOb/PgVyO+PLniVdtEQLlb5MwIL4Xyo7wtcM0Mgf1v5ae
pxAGdIHbbYvbXYEJWuk4mEGDpdLctp28kLa0NoXBbRL0H2nJjhDy0s308QvCmEOZI43qNgJNFZ/o
2P/0BY3gNtHcq1XfoA0ccREHuK++53vUZSsg5FT6T63Fd9HIndjy0xEsV61b/0Nz5MAbF/4qBL6R
47IoQ49RROvIEFMWDQBYPhKQrUI5iVO8XK0g22me/fkmpWZyxEUnuf/AEvdg5vqn2BJShHzMqiog
civOCVuKEUO8qkJ+bu1ME+V+9p9H39CQUm87airXOH4qcIY2f3yzeYpDUD1+3CwfQAJMe3tz5Qe3
8cIXqOtCzbSsG3V3ev2ZcIoT+GkynEOKicj8VPlJueIXPGPZPveZe5XOcWVlfPCzoiGL9Xl6Hoyu
u0lyfQizyQIhrGgLsmcJsh1d+Bzv2pguOYVLoACpO7noxKp0QGqb5jbunYMIdxBYiHhDJyLOh2gD
wdluTEOILJAB4sIasHvfjLbDcPRedpb+4l5eiGiKXnX7KuHkoJ4pobtwWN3iVZB1L025zeWPVlLk
sqicmT27UKyrQq20BaL7UPU0d5FN8YCNjikFV6dRfqgF+zaQ06oGPRTSRFQoTf3TRSkvAZh9+Emo
EXTVTB/4aE1aY1W65zm1jwaMHWJz6BehvNS+EX3csIcbKvhQTnpgJVDkt1OMP2AyKzejOhbjTgEH
85gOWIxL+qw9Vb4kODCa3iC2OMS4MKhNt8lI+CoJ24SJHLBqex5a8APTNmmS1AYY5e0PrEkMxTPs
zRbdqt318b67+5ef01DGmfuBmsFGhiHo0kxN4CKv19LTHxAdmy4hA9fRXIsRJiv1b4fu8I4bAlOo
1z3XJJCgbKIYCiRSxph5azI5ojXuH1tFjmZm/3buPWd/2+uRQsMpzBzLzcqmSGnEB+HdvfwwiyoB
6ktejDVUGh3jd9s6RWMaNVIrPDNT1ncnlM455QxSMJntQmokZPZW5aMouxbJWX6HEU1aHA7h1Jvx
eaU+uKS9/Q2ZpcTmIg9szA+NDRKuIubKxuOqKQ5HkfgIcep7ZSXnDOFmmGsuHSC0NLCQOlqYVVu1
KguLTFocSCHg+PhCwS2t4+oSt3+ggoScMrAmaUEMOTUzBEKa7JaLpuIkkJP5K9Zw7DUixlmxAAp/
rZZIWvfTBz4QwLebsFBDlk/yKzswNpe9YqMvZE9/ADozB2hmzhb35z/N8Ux24es9le7RjLunf923
K+0g9NFbxFTcQ75mkzAuIWa7M+KLuI9URMmtmhoMgly/wyMVOkjp8eq54clCbOVPFbOlosHCjqpb
Ji3JFnklV8O6PShK8+v+kruAXTLMKwl5/TAa1ZBwxv4Cefu7BHwSjqxcwkIC8VyiE3NpUaC+3c7D
4JS/LYoibH5w1RFZGGH0xhTQDyGCDf4JPFjhnia5u0G0kHDcs1fqcQk3Q6ZPYdmiA/GP+YDzDyeX
z2yY7lno9HmfUDHYN7+TTtIEQDM9fPwTkaNwnVAmwDIe4CxUpsBEjJ8991kObEB1hWIWuO1VvfYA
32HaQS0uzf99ZYtc6XJYIVv2+TmnLG/AWqxPFMc6h5sYQ5EFfIYlqygYI5zO8cpBBc1DUYQfrt3f
myjNVn3Bz359/tnQkq1EMISNJF9kyxibF+Phk/PojUbxlXZk3ahDg6q4qVOfGuRB+qU9caHz7ved
6CGqL4AAq2Ujf/U3nmhdhOhVtpTsNOFJ3y8ur/uQLodO7IXXM0IG/PgNHMjTBzD0wuVAiH8nH7jA
YVmnRm9I7J5fsjrVYVi1g6WF6gfU2Px7x47Knwr1F2G7NcYrsgPVyxpcBU+LMkQRkSkfN9+5iiNA
MDOI3kds43JoxHJy/kfpnZOOpiJ/aHwGvdzaOvJcPTlmf7OubsiS8SKgxiwFI3HJOOBFKEliazwR
zcZ52a2IZ/UnmeeQZBeN1m/QIV6BWYMpfuQdQMm9fS44kwOKtbzJw0OMDx7ThzI1HsKylzC7oYJd
t5oVMLpuuSSIpYwwEbxaHp17JQ2d9W2T2+bmEgR/61/HFfMXm8rzlJZiQmdWtvYznlH1yYkW/iod
SsAUv09kI8uQAQwUEtaXZOLZNDQH6yOk57U/RGCxcmz62j43kdV0ltwDTHxT8NbLUYgDW1mGdRA6
umgmjj/Uou/9bsuUMQtL+EJwCWW0/8g9nRc2iQlg0IvkfcPoTpWSJ0UxNrCQDvm4DHBMw/vIbsLI
N0i+1bU0IKdEPdmeIvBIWa6uqz6Nt7EEM8tT/oiMRWnk7wQPoMog530Y7j6XLBV69CbzaQ1QGnEI
ffJqOGLxs9GRNJ+bYnIFtZ8UTzsv7hw24ty1Bx5dKb18BKeuYOtGj3VNa9A9IsJsEFHjWei/ReEB
zXGwtL0LCazeLzLrEddVsUoxlhLdwXElLHwqx+0Ng/xeTq+LlAh7XdLER5wCcPRGWHQJ2V0aDEvK
1LZHWaI1KwTzBnmglZ0wBrywrKjK6i6e1faAoHr9Rrd+4Emw+cVw7wL83qznMEz9mkckUHVrLE0S
9HzAJ9CJjFcanQqc15VCRF7CP2lVeWtKQkyHCTxSQ92N5TqkOdpYn9bEYB7+z9/Ho1J8Hei5q4dl
DbsZ189EupJ8aUJ4h40mCT4+OxjwJmLv7GBs/1thMYGCrp4nRas2JSXspKKVzKRWq3yT2NYrxgO9
hJzfQ5x+384leC633ZQNgJwAduePzT/SHtwAXWTyI9WJ58+NHmTPDd8/+jDZkmySvrmGvj+4xMeN
bUcYHARC2sGDtZtiTb9uzu2TtqqR9pch87ULxioDJKI4us3dBFpILYYZspYnuvfVZkRqJIM/mWzZ
dmhv0PKQc4lXi0O48kZrLPtznXPW0LtF1NotP77B8uakhaSAHmKPCzwpgCI1WfOn0gXIPw+xw7oZ
JiY0O0HGUAEOnENJw+0nryFPanl5pNpauIOw24EmVG0LJC04XzBcFpb0Jdp/dzn1Qw/HA4xmjPT1
MiHLtsCrfmRMbwdYIjgtiCEIAnLJx1hmLBMLK0FvBuOmLNkXV9j3gB0LzKDNw1RcMCjQgZMxdkXt
g+uy1aenFEnFtCc4bv/d31k8UrXRjoy6aJj2j//YeFoCQnEhognVdY71tHPUl0gD2jO9PI619tVh
cXxMueDxnw8OKkQZz1vZ5s5YdlLmvtUT/KUG7pPay0wUJIU0V/8yLhse7tz9gmQMgK+mnFjAlcaB
Vc37xBgFSXYfODpbD0/NUoXwEBmvjKuV1AxprN15fd+GfuClUFz8r7jcGd5fRrFEbLqaHJfHuM2F
wA6Y4gw4RQjKY+4grNk/q3nmu9tdJel3bQRp4JwlUohROeFDSa42iWwkFhcZbSn0XCd33FnXOOhK
i5CeTbM+o/m5cyDapRPY11uFlehclhw4Taj0UovRQOM5DvUzwu38rV60qqTP0/PsyDLN7ZgGvpUP
HDlDIpqxzkOBonssjGx9usVdglXQFLhaWfc82J7hqcGqWK/OpaRTBACeDykP/VZZAy2prM/dimls
mg1LU+bHTEyqu52tI6e1GwOtqK+UxPtwUcho8xAISAYNxhxe5CyhB+WAzpWrUZL9pKREE5IzdBY+
NqjDNEbobJ/UQyYqT4Ln3FoMPbuGmFrwhN2qDGWSBPAumGiee1mu2TloDXuNucAoXeW+IFoU9jh4
5hOq+mpylyiw9WsZrmWkC9RVjw9sctjAn18vYeErpVy80fSCMzTuDVGqd/Zs2ezQJKy21H+at6pu
qB03SJ3VMTgvkvi5E3x8YmDneml06yl2yBuK0kUn5sWdsqoxjpsd8Abd8j9KuaHCHWaTd38Fy2Kr
UplFyuSIkaVR45tXH+J74iqv56QGxj3sVTxrFTtJVg3+lz5I71nWbEGFvH7sSAAPDjxSC/SRxaC3
qK9GdNqB8ndyIp4aTurUCiP9V1iqfBbujya83AcTrANfdmFvIDvcAxDziIE6JaahWbWrJxVA30ex
VYw/mBiyWrNYf6PaR7gZtL03D2pkFOb4FxjoNTZn/93AFMVa2sU3us+BiCE/9N/o1kLXTtZGGFVX
//o+eLt3XhcrMOoY3MBkwgeUCsfK0rBcHB/jqHd14KQC6kRfZrwh4KOJ8MCxgmM/JWxsIN34EIQ8
6Tt8bLK/d8+ybNb4UlaNmfBUNwmhK27HmauPA66V4Jz3cApQD6pjRO30TrwY+9bWSo1DlMxeClhn
M4GRvConsT3gxcshHn/5+elxS4knsKv/cTyEIuPm59TGHEByc2xSV5iYoVtzuRKK7URGS4rZlvyP
YFET5PCZcqtYKDv75w+MwegHrcgPayw9OAB/dMwg21IC2weBn+x4dkZQiv6fvJGsJmKLnWgZVXSX
yPAcMxVEzicpI4HMLBSsFR+Egu5FLkmHYWB8ALHnWZfh6lpC6zvzWkCnCBZ/BOIrIDVW4uMRrcWi
/8Ib2cBacA3SI1/NBzcAkksjfTAxZdEquIG5D/ZN+ZvWO8FHUd5d7D32BCfMxDlEVL4rv81G+gct
jz/fyi36yal9qUVvVN6cJIL0DXM/5S1ZAeic/UoyuzwyPkXqEW2clHFJjdLkcd3SnXt5c6osec1f
AXGDub3IibB+NZBojRacU0nyXpftiyxzPtZKlA9GFd6wfYa/T80ymmwlCjiZk6L+1Anj6t3Gu3wt
L7g0gUU3iaRoKUPjPGP+DCLC4V85IxHdGvt38UtyA3KmpFe1XMFFxXPw8Yv7lvViCpQpRIYw8wud
BoHXRB6jTIvai4od0xOh2JFWEt3WmCe152KsxLFCNu97sAasvhA/qHgcBAIv8HfrdfQoAFZAe07t
5ILb0B4ocLgTdvy3MAqfe8DIj2uVpFw0+E003LtQiRWZIjqJPNJZOLn3NjeokjMlzz2LKBZVrZu2
RmV1vDszeyX4wivRJP2TQShshvZriVkNTZL3CljT+cweM0/iqcHwqV/SqllXZ7R15AFnYiSUOGTc
qJK8zgNyLHdsVnHNDK032cGWWYsmtsNCz9ZabPilyC2XwkSnlxG8t9IekkvmlArALz3S1xDVqt2j
R+aPAIEVHfL3KVGbdZZp/YoRo1D64kCU8kd5nsEiIeVauwpheFUvmLntN2KP87KWtIhZnJoIezxF
6UTWTHByJZjtnPLzKAHVMw916RzjQruzDNSlzfXDeAtJQHsF1DBkvRU/yso4NS1xhEmeijnp4MXq
MRo+tRnVzFnlxaHSDAsfdfnk3+hpopXTAj1BEcqgnJETufpK3QofZ0rjud/HCEXd2YjF4MMbuvC9
Rbzb4QWHsZApVeZ7b8+cqLEEH9BlqTBxGmPUtbDUQTS3dghJs528RjJYM+H3iAdSpeFAocNM1/pD
MLSx0vfiU2jiReXXVvB5+ietVrKBDFqgaYQCd8rWl08HiY35tesgrmSFAYulVfXY6W5LPM5hShmZ
/rbeRz60vmNK+8ROSY96VAE0WufRz9S/meAPH9i8qlTJOdNsy7E8X1Busrn5PpiteHaemmAxZfLQ
zZJYLDZ6qhRX6kp4ZsHej6HRR4UEQAaFc0SjfEda8N43PGeSqZTJ/qOOOEuEkaZMHVK8qNgaPx9i
cG35osP60kicGt5tgTd0ZL5qytLcru5cbsSFe2YsR5rMx/tXSGcs/H6MPHUdzeFqoCESCHWn2Viy
DetY67Fru8LY5J9PV/hzsHltKJnQIcBdBI2UESrDOq1DfZWf53lJiR3J8XJyuCwsgY13uuJvajlP
U7wM7MpsYI7r/Pu24OsfmkTRTJnJGQZaCiPEA16yNRcURUgWbjPgOZ1nLNsANnLEMlpOBdAYDdjn
zAodU7qJi6s5GEhJUhlM2qXA6FbqNpNHWdZVq4LA/hhUyF3YI9oXclMSW84eWrreebEvxnY+QLlW
xsroH6zjHYuDni43Wn2vPJLxXhTHw15RFhNgxmBD2Z1kP/TLVE0T9ocIZ4u/0sJczILbZFq74pFI
65ubDRl+DqGP2MimUqjkeLpVYGiPzEQz7Bbu+aYLwn/eR/fneJVp5KPYEjJrFGre1txGzEI0fznU
8pTJKexwWBv3FWxgaN40TmRv7qYDxJZq5cdet+8IBdp+Pdks45E/MWN4HZwz9Qi30gcTWwElp34Q
gqQq/AIVCJ1vXfNnytXXKprl6dDNlyEnG91xZ2xSjfdAl2hG4os15puEeqYf/ittqaXimiYkVPok
M3nACMHVcsEix7EJomSzfJkgIb/f7XG5QH5xRjF5UJIXl9+kcwE7b255ZL8EcyKrM23/7RS0eStY
Qw4mOn6qj4aO+Oy9aL5w6zaHEwrzq5imMQ/aqZ/jXhqCHvg8WQuFht5plLIUtoLdaMPvh64rbY6f
JypnGSf2M8/iaUSrw1APBEBecZ2NaYBGoy6ayfoQh5ZdVLoex3KngMZDlE4ZqKeqLDhUbX4TMeCJ
5SQvAERHb9G/RE6ENArrWJO1vMvGpxkp5JeBDfAKDJNDE1pTDaDkrUd20P4LQEtXsckUCJFCNcVn
7hfEs11wq7X9q37xFyaSPEI/079GgqY1DuNSsq254NIni95XX4tkCAfvOdhiv+Yjx0HJIX5waR06
7gz6yBqMNu5gcp8hwjgrZiIxKUQZ7lCdgI9+ZeqjVqo1XT+LbMsCOVsz3eyIKvdlcPEFWEo871P1
A4SUR5Q1wErkf7vz+pa7rxDrJ1A9/i59ZLuwnfprRbYFHT4xGaC0amOWnpBYWidiUIDyDzCHpRsz
DFGGylAYW1L474pzyp0CHIaKBruEHe0RucyFbqJvTXbIojXauqqZ4eHCmkCPl1incqQRC47MGEZC
JIkaUafgqJC+zxhOcpywu5fgOJoyjJl1QpNEuMmre7Vq1KFHtdHR0yoHfOY5IIkIMrOGgEwM85cC
mbFN551MMl8Stwk8rZWJ3t/pOIyiwjk3V1PvNG9HrrZi4FJ+BPGtzq4POSxlSq/+iw40yqgTG+XP
DvMT1NNpyXe+HVOvnyC/wpYNp0RDZO/UYHVub4DGBnzWtu592enPhtqqFaGAeVxdC38uR1FjuVFP
VZV3HYI1ZGIHSO02IBxfuT9RV5VJf7HsnDUjzQylagp3k1elYkBX28w5b+iXvw8LjpgY33b3oOrp
TqRl5aLrUVcv6blu8co7gGn8Ql7o2onDlXQFvBA+14yQgBE0cccJlBDuH8YAiiK6rQkcEYVJ4ihx
BbdoDLPKfX8viNgMiAoFrznd7iJYgooOB9X92gIwnT80T8BASHIm12FV9k0yuxJTA4jvyFDA2oMw
uDskc18JzzFANg8cExKQBEFBMBzyK38WywYG1bzZe6Hv429u0qdCEYAvCUl8TqZ5sKvn9LxiOoZM
hTFayDZoLysY6kXc7VRVTyG9K5THycajZHQyV65v6Hq8fd0v5v3/W9yMXKXjN0k4b77nAN2QuusU
/D7C3zvP1xiOGwCMGBjN+680iH78pdROlIJCFkkEEGQOUGrhGLFEvdxrueJxLG7B4ZuZXw7A5Ich
50EAwRMuiwG5vxYbVZYGWsid8YLu9j18448VYis7djb5tPDSuBlqKhS3qzN94YLjjI7g5Ss9bOSu
+38GoDrATF5OswdA6YgrShhZVI7LyK6K5ptbf/ofdACv4QJ9ItP4w1tR6mgLeIhdJi96BErDNvaD
sXXIipT/7l/yrByLrx3K8DmBGbcTGM3VvOdnJRsWoLnLNvpmZvPIRYCai8Dugj46m0uKf806i0vD
8Yqe6BJVRGDuS1otoU7nS7G9y4CP2/ikAVeuynI3okTMgKK0FcM/nmTLdqKtySvXql0VxrLKwBiF
MHzu/NZM8Fa0YZSQpURsgQf1HX+SQ6b4lGhaG7sDFhyeNnbV1KU3D3K4dng+UWPg4sheK3QTtew1
Vktw0R5+74J4GM1l6NijUjLzwn6DHy9Gf93DtXgJHR0TFswWwb/Z7zm0tUWCBaktadbviGJ3JpXU
6fvTL3Cvny52QDIqDD6YxKHenUYRN2qCfxE2S0H9i1aVkOOjLmOBTj5jut1hvT9wXs+HjMjyKsnN
/dlKBe/aYnXDXzdWPGOYqDO6cGKO6MKUxbuhhZAXKCc7wurf6neQfRLrBonPqCIliK/Va2YLmyhy
Lk94n/o0kCT47MqguFBeRi9O2DcX15vCzlS6ixaZkoui5lsUnddfrvrI5X+G8EcwcPW+UX/12ZXO
I5i1C8Z/OT589eSahbp2HI6Sd4GqfYaHqk8wzHekN/E0ZTvSxfKHwOrbF3EAd1JMQSqckpci7kpU
jqYFy7bDFPSqIDw/iJ9yA6EqIiS9lT8sIW5mbNTeMH0TYdy3c7RZaX8/r1WgQZhQuWwCjPnea7HY
CxPRVAblZ63CzDT9Tjx1GT1NAmgTr7w217NUWUG51l6RlMVsxmhQScJUgYSm3+gngTfRCeRqLwqR
ulb4zaBcJxK9TWzqrGx5q7YwpfWbHTDa52JBkV04L2USxa90tIoWbrp4QvyuV4u4joPUaNTOy/D4
QY3xt4TlrsW8h/OHB2yty2eTkuUR/ghPiT95RrnzkY2JKAXIwLwr0bzE9J5oT2UzoXna0n/WOlCR
0vJlep17Woe66guVz7WINZrJw2BgBOBM4DeUne5T3dlgRYKMg9AO4uFpe8KMe02BRfkBKkhAUH4G
+EB9AC+/D5Wl0ghaUA/MNTsmh+FlL6JN60BgC4fOPvlyK5XBCUUoek4EEERwiw0W035cfTsdOmK7
smHNeH+FH9F1IAtqD54TMacTjsdf1Jou0rhlgSbqoWH8q+u0njglJP6338rvi12So6ALX+WUuBcF
CBXDRfnbh6t5DyTjrLkzgud6EWdqarZ9993qDumB8TR2Up8A/O1B7hGkMU2428Da6XLvezzTLCte
AbBfmjZzcXYoU4KVZt6/4bpX0O+W1Wy1cdNjtRFuH6ndOqHwnXDXYLPtVsSdvKoZ5Hl9l1RegtqY
+r2t2T8IBRvNFvvy2W+th/x2k9siRD83QSa1oghnxLVi0ry/tIOF+GSib0A0d7d3JW0fSj+q/i/h
RbnfiK7tH5zxa6GLn9VjRNWyIlkCp80kiEp2OcqedptTwyVgmAAa9g8k+UJN1pzt2tqLb7wJWKDG
gZzU1Su4IvzeZxkNQOZi9t5CJzJBdhNWBM9XDG9YKGuHz54ShQLx1MYaP6eTH4LMi0w7yiMuWt7N
vXpChutEC7swHp9FIaySpkY1BQOyI6OauKNCyyngSudU/Q45L5Xtu1WlHiUFJLqeNE0zi0tJh6wN
F7PlAkxdEtoLVcbCe8U/+7wgMVCWnljz6w6vu2QSvRPJ68X83rUiUwO0Z820kIIgUeK6AvswSam3
QzRqkUL4XaElROq3vz67d+dCvyVcKJv3qbQqr+UDpJnqtoyL3/6Yy7ijAuMzyWCHzDDf9uHD8DYw
Fw7qFnoKFFzsxy0FJttUJFYDR9lAZEOLFGbIKtkMG6FyJF3RDFm+dwbUj3kZ6ge1Vk0KxiKp7dl6
QFZhZ9LE9zKnBufxSLs+hpTM3tRTu/ZrOX/EHXRw6cAkl3gy/YAI9Oi45m0EiYud+08TWLipDfew
SfRsbIUxB5peegShf/iTeztBVr75F2Iem6qFGBH9oxKlBKi//pkfcZVEeJKr8TLE/e7BSkTUT88N
WHp5W8tY5S8Z4OiX+lSxoxzdTHyYwFYuNh7/IOYX2pqZGNHkNCpY+ZAaynoV68WygEOcSdTVXLu8
cTYbY+6BdW3MRVQJOitvApcX4VPup8lKYmPqL/F3eS2hhn3W91GlbFi3Nom0W+D32e5WC2IltB/5
f1Zsj6uClMkPaYLXtMTf8jVOztXdOO+tDmfZuJBwU68m4hQmLnyq9WWNOw8lqklS72KdUC2V7/cB
7ok0C3ruqlXKDcv1c5FtoVkiMEkxwaRjDG4iTai8GIJCvwVg0McjViW6+O/ZLW3igUNXC36oWKYy
ATLeu3eJGe4bbcyBBJY0ULVih+q81hcwd/MoLw5ooJ6CgHRrGgmcC9lS6/+1EwRiQ2GpMrCouUVe
Q1eUn2KSX29l4IcIqcpZxoIrJ0zScFH2UVIaQfJCzSVUCbx5IuMbHQWjFqD14Ixrrbnjj46+E3vX
BgjgdH98wFbWBc+TGdJHU0nwbyI7uDc/ic6QmUL82a0N5m0vr91w4XobQuMbrPn+CM6NcEQWk47j
mgx0fpdO94iq/RZNJBS61stRB7/RU1SmwIBrZRhKaeiacAtc8I2CCW4q33qDMsgLxEl23SMzuN2k
BkIiZri/jxoAsM0VS7BA3CQ+HhybHr2iV95zmS/YVPNEMu6O1CuPHchGDivRuai9CWcGyFd3cmZ6
b0sPDYrI2qWwkxqhIqYljs1TPNJvxJOJAb3ao6DWeW5oPOVtiSzAnT9E0jkwzGNJWclOHWs6Sf23
mm38AcVxhX/NyTYG26czJNBw6yJIay2UqabllWrYRGpcrk2aekjy2tDWLJjlLdW6kubuMikSOWc/
CpyvC6VLwB7pJcgOa2zwaUVIcj/I8os2RRFJ2FsCLMO8M15lF3iqO56uoBuHgYiG2FoUM6lssy3t
A8DIlYm4UOH868u9y48NCYuptXTMt9h1l5909Z2FN2/tCXJGSlC600oQsYVdWSNO6H3na5iUlGo+
WlUA1P4GotV8g+W9mNRM7/VMkB38+//qHN4DiJ/YT295zJDiqi85HBU7bsoDeRSxJ495TJfmUT00
pSjDCo5G22kGVCdBoQ2IA/tOjSZrteNMiIbJ46aSckbiwOOzNuQWOW6+Pa7OKpoyZMf3/ea9Zwzx
kBBAZMxRnWHpJBYftvetBSnrMaMTi1yOGR1WWjb2/oCqXi1LguUik+hsj0d9ssCLuOfd72xAoZ2L
0y5Cx0r03beIAHdyJVFxzN7BWIL/7ozwebz0szAgTapy2YSoCNpCV3QiaBYglhMzILn7fCkWbNpg
QkIeggBrfFE6Ky/JYkIsdUHNZoMALrGUP+o7pzSmsBtbMslWmaDUGhcmKMPYWebYY5hm236CYjMH
e8vzfo2QecPuKb4x63O+RRywZUaNHyIW2cxJrcYZiIoiyMZ9fAq3Ze16AqfxEzKmu4FFjVPY18zp
Ngk1mwF5jhFX5/wSzByCb9SxxTGamnijo3s2cR6zBA6aqn1sIEz+vZA2HrOI4uqcYXKBgQyuXIOc
rJsB4BA7p8/SgoSBxxjMmq3Vjje3WrnNU3UOEdq5A5XSzMUvNsWGoB/PZcyeQtxD49f+3hlgsvUa
ag5jzP4+ZqZXy/QIG2fHTsRE6oXKNatJKN3BZbICj42nM7dHKzd+hRnvwwSUERoVQoXnMmXM4n8f
+s9rKQo+RkwTsFijJTGix9F0rGTiVI2qIQGBBTakKrtgorDCB1S0gI9AxPBBUOaM4uE7t1RdnQ8z
cYjcWt29apy5DeVYupVVc3QTOrBctme5jebguZvausJ7zuZ0DnLGtK7P+I5n9i8/AMCWaLMNIQNy
molQIzZ3t5cRTyg4LMS2JSBPf8TBGUjRqQ1jE5NsrUzp/ok4sHUfIJNA1qqbb6Gwpv3XhnWJDuBB
SptAKPiFOgzIinbM6af80nPpZdkyXd6v0K3cBCKbVi8uwSbiCmzF1guh3I8UPAzI89+KJW7MSuTM
3lADfMx7+W4HymtTX0XzSCrf+5/3efazLxx3xmC7rnaFnzvlEXe0NztFmC67+E1kvPW6bFTlbNqb
HGX3uFlOjHZvD96/bXCc+Dgjdq8iSxCUx45Ut7hGiXP6Pne/4c8T72avDc8nbS+eJm8S2yjEdw9X
zY9gDIJVFmVGU/1hrcObOStS1S1v37VsTVj23Ea5GPSfGU9M2WCcuteAXEVsStrgBxNJegdriEMy
eO5g/KFKuEmRu67szQrvnRfc9Rkq5hh0X28dCmbrOOem+ClNQYcVINHScz0IIT3Fe7Thp0DNJGM7
MWxR3qpsogpNGo0WzqL3dPRr1K06nabhHWIaoEBHJMmvv2Vf5Ai2joq3Ne+vLN88aZ+CKGNGI0Fo
k8xYeBQh/C6U6x1mNlOOdMB2CNAB+iv5u2BCc3QKYFRMzWby5AJ80hvpHCfcFcORibCKtCKW3BMZ
TKq3jLIv/giCqwDsuMxyfIBXCfo66hoCeVTMsww+Jym0hSziNyXsUeJnrZOgN0fJ0oN4c99p6cin
5fNv4L4wLTVhJrtLFqLcbghmy4iyeYkOnc2U7ruUOnUWXs9oUdPEC/N37DyWiTUDP69VkswzUNmk
j68lhBHwsyJH3O7FWH1tgVXl1YQWzL5DDl+3nfNPCx0ZVdH/xN3ARTHvVZ7VU4DXp49l4O2DR4Wd
dlq8jKMmwIn4cYelmMTPa0/WnFZQBg47DOwgxDpuIFt0Ds+uG7SouIzkbJSEdcMrLB16vPvI5Z3Y
QgT6CWbVNd733AaBbMRl4DFenaC80kkDZAINoq4aGSRQ24OYCfofUmU1QWSPw9Pr2TJWfLexvbox
6FJzsgoqJaMjym7mWyOA2Z0ZAQLBhHXIcBBCawzDp02p8vI8Sh6ZqHLhWfA88BUwlW62VMpZfavt
wmDLDWXmwyK/p00wto1qxNBKVuRUcJsRLf658CIWmDJKYQWQ0QfTJhVWd+noNjlaRBYjSZWUtNBv
wztfB3Zv8rE1k+l4wbSp5wSSt7ZvELXw+rRV4aVVoERJofLA0TPReE+3yiHm127J7RWCF7BRVW+B
h7yLj6Du3kvjmzyWhxOZV05WdzCip9OHrbI/5MlN2wvlUEdxjlgH5NmL0EJ/xHZvc10vcgcJf205
10HVhrs/Je9atlUwL11bLBatXu+WDsK2XBHa+E4CEffJl6UDGqu9aDXLovwk2O9vy9a30VZImyu2
YWoTT6Kt0NG3i+dB/4L4SFUtOlAaSzThwwVqnJCu5CvaW+Y2h46+MdSbpn+NeE895ReyPuvI55Ib
JL/FisKIpLVl6y6jcq4s5KzN6yrxisGqZBiSAyhcWY4fvUbQkox5e/VA8uglWLVOPPcWlLaFI7oQ
gPkqnAdtha1ZXFP+mYwQWoVT1WD6lpFaK+a3sBILyRh4gnfZFSvR/aAOQkEvEth2UJFwk8s4L1g3
izkhD9s6MY8c2bQTuaDagdOY/uwSwanJ76Rwg9HzltPuaeTmMb1IObZKWliDUQUDALBWueZrZdpB
p79iGrQ5KPG2gFGLmc8AMVkSGWWPcpSgLkOyVEmPGTY4fAf7cyqaIdK1o1GYQqmzixMWyj5X2DBp
TNE0l49cW1guAOcVcGqlEpN0YSepmo911v9JjxoUPiX6QXMajE8nnloU2fGyS+12Dc5QIecn8eGB
58zoV4ZbBn8dlsVAoJj5k2VViR81yleGoiDDC8aZtOi63QzlaU9WS8Q/dnsbgmn1MdBEvwmrkjfr
G4P5KoFcF0PuvjsdqTq7uSTVhAqYpCBnhQBHGir+vzVJOJ+Oazo4FTizDLn/pbgI+gmHYD7kUi45
uVVtt7DJMom4pqw6pIfVCF600RvXOe4PRn7yiTBLgWbSull8qkBcl8DSbMOymPkMtif9x39lKG1r
BdjpT0WazxijXTEBTSXZiKUkxuAqbq0/qDJlsLy5Kyl2QwgSJPMxsxzY/Qqhtb6sTivg0ieFas1n
9/r7wwxm+ptWvGiUaLEa6Ns3LCAR3u0fu6FtPf2FZw/hnNJoMx/qEHxGG3XzM6pkayq93guPB9OS
9hPl95jCwmPmfkjziZY53ZAaUIKAkb+gGBCASr6XL2n6R1zk0j3zRZjN085o+Oq/9VzbtimMHgVm
uGpNvUHUThU7Go6OqnqD4UzhPb5HgH9PGJt+clXQ0a3DOkl5KfqQPpLd/njWwb6tPAf1UFyW0uaa
tsnES8KPTiGvXlmASZhY/KJ9qiZIQU3T7gBBK71eHPne1LNnjq1xIZi0oY1ZvcUn2bo4HDpTsHTg
yi8x00QfkJYpmwclkbKLVINV2j9AJTMQ7bwK1f7qdN9OLURLb8+ibYuPEJfFOQd6DPJrEIQHTR3l
3FSXfLa4P2nujb3pQi+Mx8UxUmwl8nnyufQxFqZpxfz2dxY9DQ4tVv9DPAUcB1+/1XYnQrCgifs6
qRcZexMFVxcZAhMabEFxZVzA+oedTyiGDiMqkE3DoVmrzIRDlbcRUZESQ6U9Mt/ZLSZ609hKWHHe
b4gGQEuMmIUmeKREcftOD58OvJDpGRcuxaGh+HFIXv5qs7KAu6jSYxHdjkGRKH1MrRkAHJzj4oWv
9swq/xV0gf3nFIUHyg2MM9EYHnryr42wNtEtYzfDAz1YbKkM9cWfcbHQhPQ3+0CSkIQ2IMSmr8JJ
VEDDtBi0+xuE4jqco9j+/Lli0VV4EAZh+lzQKXcxvGTfPQ3wXq95PNPHIjeFJRXqmlGtE2MEh/UP
hADvYBYheain4bA+bh/2wFhKFUDtZMGahpG46jI7Mn7Ii7DAVisuD1q4sXRSoRk2uMXiLtvY/wgI
J7PtdT6bMTAShMTWi/CnwhOrcrunUX58OtsEQtAna/+4y2H94exFTIkqi8KxBA29FjEagzsWniiH
THwKVBE1ecZDGDZJOeUnGjPEePBNXlncKV3T/0Sbln92Qz1MdEu6inxrHD9Reb6VTXpuZhwW/up9
hmcvF91eFC2G439op4m4IZa9y/V+r8s9p8Qi+73mjnYwvNPyxWhtDvRJZLoJJUJt36+rERe92Nby
1d8bjNVD7MXDR5SElCTBJMV2woFhMGyC6azchffb8aKFB5btGB9scpRhGXoiSajVEQWP2aQLGv+r
RsONgyEX2BuYkPydeLdK0SLFpZ8XAOZHn9Fw93BSwXLgLuPG153DechnwTfDMWtPV1SiygwE5T0M
45QDVlsPc8lH4uRzGWcc4uTFrRMmeFK/edVN4NMzOV0cdYXYrAO8PI9xwDSOpFzpfVqYyWsRR4Be
c3b34x2bIwPblKZQ/a7aQauzt7g/cSZA88LYSCdWiNjOsWmIFN87kwITew9oLuHMNfPkoW2G5kqY
7F5YkjpPSXnpIZDhwj7sef1Y+rkLQ1WPnzEvmdUXzwuNjFHSLxGOzteBd799S4yPR+fHVBTduYkK
s15uybsWGguSPaPMS+b/tf6COVCJrjl7yHvwoes5Ox2AFwo46ScfCRLqC/eFf1OUvK+rOf18OD/H
nNInQDGH5gwXVDR82cl5O8vEID79I9Vu/ZawlXIAvZ5x9MCnPECSCgk6WyI+tGZ5+XmujNeLdH04
qC8cH75j39S24qL01eY5n58EYoI1HMAaYgOWaUmCAaC8zva0Je5ngQ/A0wwl1Ho0aw0PSAfSYqbJ
7utSksG9oi4iqNEDPOLruQxRme/xnSE3w9StH8BU824t3xoPRUvXhTH3TQ/cEwL8RIpU+zHKr9ZM
poi28zfSXmLZF/FII5Hu1+NvxQgVz5aIKVB/AYRpFfNIC6DmRkGMobRzaKxMQwEbyJtZekyoDzcU
9wWxXlxD3Jl5cscLc+LL9wLhicJQqM0JDE/RhR4tZ7COn2WU4e487Yfd06n2Env2PrwkWJgRg0q1
Y4CV2YQjeoaXxzXaXjTgLHVkAm9OeTzDb+CmJkPpTSI9RmjxsnQO9zdKBq9Ilid6+CVxa8E7kjVP
ApxBbhdjNmiZnB4v1e/q0kJ6RP5iMDegiRJgpJW2VW7F4jahd7+s4FQPDdlXHb8X3tMFKylvJPPU
MHVvAYUlQV+mYV7X4bjo932QuBgFBWBEJD+16I6VAfLOQMxIePtuUy+C9LuoOOUzzE00JNaDjF5r
oOJYwP+3liwpDbMnIeUmQAs8SToW/7PwKKGOqAyVD9Wq3w+0eaD7nCYGUogsdMUqzrPwbIPx93/F
xxtS4k8C9npKDhwcveCnUIXXQEJsQ7tZqLbN/8uZ3o1wayTEP+SPd3uYK524ILNLqd3EkKNhaIFQ
gYelTIO6JwTMWvsHpqU2c7CNLzhqJaoNQCp+p7DtDpT1Qe94y0oWyUrGLYZTxBhQESTqMKcX51LY
mYf3L6VztvAgIQ1PpSH73NbcBQXrNHrN7OfFvWINwpWELFCxZL2+gRuy25yhRkHT6Dru6KZNZ+eA
cPHol2SdhfdT+i/fQZWzR5e8G7EIyL8mue8VcbU464e3ukXS6gcKkAWSLJvmvf++bq3cVgc56RkJ
SNZoBiGe79TuSyUUPwRKL9A9CYInqZGuwqqqelebMxLCluSzMNLIzjBR2WaIcTJjOUTSpjjJUmJ7
Cc/XYARJvpzZWpkbFa9bb039PlVkdFz0xarSgPFq5pHzp6aWDTyCqxjeXAKXYp6bcNJvHZqxLhev
WhGqknuo6YTvxUIv9C5dFORJRkU1dU+4l+LDLBCtK6bOmjluxomGycnPrXKk8VAPAJNdLpL5q/0G
kFH8iv5uwVr5BJmTNXBjKdTudcuHRtfyqsbg/1AOoOfKtyHPs+iDOA7c5oNsRo4m8EajTzFKMsPi
Hd2KraIyrqzMJdHr+VRy3OCDQ+HO6UFCKS6LCcnPS1+wgXsg4mg5tgBw/ArMixYvDFFoPvrWNnGR
duhJFPNZ+bLxDRNUAQuDKqAJHP/ROHoi/FqH6Pok95fGbenyr7VRARiOgFjrFsistooiUVn3dj4n
vWPkQ6ne1UsKcswcUhmqRbNh7xxgHmkaSY2wuxH0txV+dGHEdO5yOX52V1dq6MXeQdEhtAaOrKGj
F4LfQAuljLln3jsj/iBaDwYfDyI4HTrfxyHr/R+hLJUkqLMboOF9KzrGiJyvLngbaxJclaqqkeX8
0kGIgoU1dSL3Yx+P73WnGgqb0SkKJQ05WdMpssF3H8RV1XV+k1Ify4yBhiBG+qbod5dQcoNcCcP0
uaGbX8KE528BaI5S6NgnnV1VlxJIoWIaliSh/5992rqONv4F1Eqv6vQ1Wer+MhT7ZQWfhRiEO83p
dtE89vK6Yxlb/MPem7vxunnkAP9KA6f53vhoZuCwuq4th+IR3TPExdMxLO5NoZ3n3uHxVJHptNaH
kpn1KH53YodAyCHUYWUye9aMjF94xpJinbjYaB2+J5ACc6rCZLqTB0SijE63hSgsZvrLBsfqdiE3
c/ojvOg9zxK7izFviWVZGW5aqkKoJ/EOzzyykaIXQ6TSVHgRVFlU1ASEovvOvnATMFkwpwnrZ/Ql
6mnhl6Vt6oxXR0FmoKNd11iwUo2xJvmZYK5cvnywsRIEejwBWoepbMQWkhVTwFCiRUPDl3TfEN7Q
rDzcw+EGtne6N88pv2JP8IHkhIdGqBBw4ZgAEud9HEtOHjPJ4Qbxiso3HMyG2LdbuN3PMiNkOeTD
Gpdukn0DSA8JgHnMqsIBDMUa098vI8QrwYofT1nJGdRxXlr90RpFExf1evMiW2IuvyK3qaj8yh8f
9fG6n5Rf1BgtxjBkLs1Unr7rOP9Tak6a1nSbmUZy2d8I/tu9UJ4mWSoCSYyt2nQKBxb1+PxFqJmc
NX5LOIpLomoxeFRLrFdF8E2Z6sRabfP0FsYVPwW90gbPomVJaXodPd00xtzkHWQoNofhn5EhatZ+
eHBpQHI7D4PkEWdMYmRLrQvDeDlr7gUqb9yG8rpFd1Yye4GMYFdoJFgkWZg1F0ZY5yAENIDL2q7E
1RJDQWfCfMDBvJq6HfmhHs2CTuYIbsGvrjz0xxDHu6C2fi1CbPt0OOLkotmKAQ442MAzBwt+BzLu
22QYwlDTVwkKDDHH6eKeLlB2Fp+BYJlUXQ+k5I4+V7O6obxzy+zlQKxXLYQk9VnxnyjZn3BAZcbP
mSLoTFgQwOwwZhUQ+8O7tWnHRl2RtYzr1yOYm/ldakDv47Ts+RAIshCFM64Zpca+m1FJXJyQH3FW
02YV4faB14wlQ1nKtfooAYLKfSvATEoJr2rsRtte9Qr2dX8T1YzK/YoA/P7UUGMybw8Ri09/anw3
7YpkoDNyGlri7ZkLzyg5+Qe6uPZ0/X/QxYaKX91FT+sTCtoejDIflPfNWLM3KSh1efuMCg9pyGp7
db1IDxsbFfm6iNbMFfjeyzYnQZsm+2ypDFT8GI2OPVs7rnltO7iPPq0lv0gm2ICVTkqb4B8FKQDF
jYHWK1Wl/hA5UgRw7S1wJRZ2V++GWpe6hS69trHrtA7rUJNGkcF6V1DWYvRyLBKf0HyirxmAeQ8U
3VdoGgXlqLBSN/txVx6v7K34lawYPO7snEzZSCnedeS5J/Rn6DG59r+E5/KkjLhzAZJNulBZqdXn
9Jy3COsZURpcBN1rDbfrnd9A9Nk3Ki1r/phDd6ukUnvKWV+UySxoJVtbr83Siguf8EUU+rJw4f1F
zz6RazPp2SvjL3EEFEhZ3YwcGE9zAgSMTR24ATjm2bPwOJrQCiqXhmKgNkYGl/1ORDzpmqqb6a4P
Uam1E1ZmQiHwf3bUGkT+bedFUUxGJ2ghEt6aD0pjnj2hZMLsVZYpiLXWiUagHoYgM4o5F8+0PzFT
nfRhGfst4EDAgRgENoxy9+zNWpyrs928QGl+QyeuYsXEAx5KdFsOMskqziBmxVRZIBv9DGyS6uvl
1AlS+A3oc368QKewa1NFRsVf/0CwyJVSGp0oRf3uRppR/rQSkO2YUnz+jcJA/yTX+Y5Po69HKxeD
NLd5ZGNdXun86B8E9MrVuUiXLPbQrunyrtIGhO/WHjeMgoTi7NrrtnjzaguQc7WWwI2VHIMBam32
UrMonfIP5Dz7MrIXVWjvT5xT0jyXtu1Mk/6KkMF5x/9WEEcuAAgJ9erRr0c5bzqfxQ2B1OCUeAWU
l0UkJStYJX8Q/mrJaXehKTKS7fCNUT73tPAqq6LO/20TFFTtTqLyhCiKJl9c45vUZVTh9aoh1taJ
teZ8Q0Y/r2E+3ddQ1Nm6+Z0BM92XvkEX8yhmfpAXFpKO6d+8IWDJvxntNf38Xina7plLUykLTlrZ
n4PAHilI0zMBR9aKV0YYvnwbVaOi3dw/uBBbVfc90UasmlFT9nf7jzX4NAKhq7gbK4UAtcmC7ThD
uJGWhJZVqIIOJ4FJAHZLSkCu5Z148qxQqyatUzCkHrfOQuoBqNQwvrLMUmvdxsBi+yiiqxt0WcXQ
o+xhh7vkMELqUC5GXXJn/mstWbl12wiyJxH/EIcE2ZLs0KzPLFv4ZccK9y0ZqAvm/lHRyWM/Yq+Q
wNOTaBocEpyu08CaudiiEUESlmkYKIntN9a3AwwNvENhZL3KdTEK/2d/Dsn4PUoUGfEnG4xZ+NU8
dqcYiJHC1RJUHOb7ybvmutFfsgg7OrqxvS5rprBUTPDEQjOLDeHrQ2JgnStQFyecnSADKJrP+xtN
qYi7srHZXflN665l31IO1Blf4UTgyPRcwOLrsdboZd+He28NTLWHJpTAL9RWgCXMFoiU8prFo/pi
w9BeVyhcsdMRTy7+RhCTEFCJQtMmVS0zy/NpwdVeOMD1jmxjTajXEOdOJDaoYWGuAj3TCd+jAZpj
nFViiYhUE2yh2MmuP+TworLFSHx/xvHacEf2ZyVT+qcI/7rLOsiE77qjdsIh43HiFa21rN5UgHM1
AzC2/ZvjrmkZ+H8uojR1+b2ofGj9TKYN8CUz/4NAsYoT/F4tjHdPqeNCEFqPhKVslOfkgoJ5eM8W
yMi9fbttPQiCoAkacLV2u1okel8jAZ1Tu9Fuueonn0DRq/DrRtIoVSLRSi82wwUHQ5kh70GizAJl
AucsQF+YptfyDKGafdAi/EDOLz++2DEQHsJrYInIBD72kT3hiY/40zFuDFcMSL01MzLAQ3aChF0n
J6Dk+/9rBm5bP1VtE4BEo4M9w45cXc9aXliT7FVl653e6RF1PlbOtBOgOhTfyFUFkU/R+XfCnwvq
6fVxTOS2aUw0guYXZL+zAXWmx1Jo3V2sv8lcB5547OGmPwbaL1ALkP+3N2d17plZjYMIEz2FqOCk
kNlLskwBe9mqD5kuGUEQwbjD++LzQbSajXc0Z1CwWGipUJvnCSlJLTKu6FO+wiQg5T2GfmnjY6F9
eKehHHg6ZyOx4iWXR214VTKJ8VktV9Yizzv1enMc2XbEXvZjxaC+sVgoVdrwai61ZVukdYynCFPN
8qv6Acd1H8MRTt98J9WiQuWHNDREkg/BxrR1qaRK2kwjB5ygSO5kJEI+kKxC5pS91MOkUwO6DHWc
vhRXrKBABc/49rgOWokiM3ejhjwzsFBSxh6/azoN7FTa9J/J9YYY3LQHkvfNiUdkRIdnVFWbU226
g4UjUL0MNKUr2KTHfFRGL+iD2yowmLbLcYPUH5ZlEwi0/hJYMb4EtDPzLc/sMGfXBdxeTtNwrREJ
OORYm3WnCKQtafX1BlVrG5xtFOgE6aAH9qmAJBFUlPjGZDFGXhew7kDxjTTR2LHoQEcckbm5dYMc
v3kFBxPoiZLqY1GT/KyaF6XJ0w/bojErl3jLvMEfFSGLYtUOgjzdJjPFkZYD5VOJy292jEDvRqlo
4vynG0EXmSoMXTTpSjhf5rSrhQ6VdKUFh+6wO8nzh2RPlreJIQjxbBKp1R3syXrbTZP80+BuN1eN
kSyd943QmYMRBlbrd6eZD2eDmoK8FWe07VRO7GCnnmwn51upLLQBW0b1X+DFEigxsS4kUj3JOQVI
yr+vIK23oCyhdUmtD1wPTQPDx31nslXChBVnBU6lX4OLvAKY18vr2eDJ/IZHVRcJ+HEi7L3AmkJk
jqzTScUiaAX84dPJItnHLtgXHjSlbGdJrjtZYrF8vcncuwWM0W6eIx15psxijQ4YMJnJMsTqZQrO
+yXazi82J0x/2SsWCnWMwS7lsHsPrrHMfbPWOOLaU9YRP10bo9pTDf/xU8l+28EwF44liNATX7Bi
hExSKbQPbi8I+hcltYk5aE7t45rE5CsoG+qGM4pK3qbiPbeksYgio/kzq9uQvl5LC2RY9Wu+T8fk
l7zJ+OZzul9GugD015zyXb8kpZQAtijAx+YQUAJqjJLw5afxYjqWeSiWMAA74gJ74Zs0defUB8Z9
UxCN8Z6pZE8fRELoO+R4jgcP9c6FIFa3tInHVFHLqdCkkbcVFlawenN22+JWMcSKFqlxKMS229+Q
sq44C7KIaWRgCquhnbBwKSJL+k08dPOjt+5WR5R0Uy7OmjR4BYLDZPlMONnjwpkp25u4gDsqqHIq
c+DQRhOEMOkf2NnjJAbB1vuMkFNSfZ9j6ESu4HQWd1iCzqNsHI3dKUpgKS809gIY9bMZFwh4Hg7W
GULIbpYM8o9JqExn6hBbdCRAIzC4OimR03Lt/zCLU+BFFWeYIgS59TD9Y2d6vwvTpr+CNqcToxAX
TUHtnt3LCgqspfvVpPvoTNXaS9jLuEfs915t6LCggJ3uWM927R1bad4CQVcomIGWpXh0UMRs7jgQ
YDKP7fIgZcNr9thDi1eoOTipcndO4tBE8scExUQWwxsaYd4QhpgXYzl2OfbUj5bXBL3ec6H0c/Ww
7xGQcdBAwBcE8JRp25hxTbVoPpIYUAmrP/g5u+68vnHb+LHRqzhSc/ZMpZvnSUQ+/B3GEw/YcRTw
mW/0z2pIMEYj+Bi05rRVfRFAmFK3Y2ef/gns0aUYvLEM0krDil6cCPlcPsdlFDohs1n4hhMrbA27
SaRkT/6UXMnV5PFkYqoj/fELj6BQweGLlX38uOfObSBzCsl3DH+Cdg12M9WplqQwhW/TNxpfso8i
wVn0tYQWJoE89IsRjJxkAiiPG/WqDY4CKV800sYAb54l81jgjrAemilqlOdk/Qchmr9AVmTuIedW
h/wxnPIXb1XbWSPh8ddFhHgi5AJs97rBF9Ki2HsgIxEmdygMX+VZEEjyxYZbL+gMhZx+nYhjy8MZ
KnkuRH1bq56J15a/Ndsz6OL5bfXPVfTG0s9/m8o9wCidNN8Av17/5qwTffxMgxMt8Tfhynfm4GuP
ZsgWTBILTdOFimt2uMpJ+RdflNWRPR0hMgHRK20DgAFd49c0EucdJPyprMLxe7fha4ZT6oHkaKLf
WBXPGb3HHx5ByUh/5um9RWYUKsVGIdcLzaJ1PREMjYA1VjilcOMA+C4B9R88jQJsCsggU0MphlLu
5BdnLIc0hSExu6PhbDxOg99+i6o2cA8/SG0zF4ZqUdigG+6IwmECneanYwdtGIAeWC6hMvwcSh3H
rE/+9UT2p/4kfaTaLcS0RLmK5WSrfNCjonLzcYoJIF2UAI8TMXE3ZXqgXt9HLbPx73cXYWNrZylp
TM0kfekimGGQxPtMLrpf9o4lZVr4ayp88SZ+n4NL51PR2maeEpSyt3Z254Bsh/Hz5zVYNs4ftfR3
7Zp8/mvsUl4RtYLOm0n1b9CUGCftx9xQi2fLNuQ3du23miqq7XRb7hwyk/WZB3hLXrOfLp4d+6mt
YVDY8/bmqnSXi+TZUezoAv1+jQim2KTp/sNsq9PtFMmByHzVa7sCqw2PUwHA09I+dkQXX/6GkWXe
/17ehfvEPtQym4NP1C28E0fMQnAhub6SLWp2cpxbNaq/zuhJBj3wa6EwgR6mnL1lDgCWW/Ubidcj
usS2lWLnzkmjTrDz7ZnydJiVZDrGoSzXV5anJqPNrW3zDOpSrsN58xGB3rQbpUrQSyl5hN4nn7Mw
LDot7W692blPkamkkE9wG6PoMBlfSopalnKHZDTtduPoc7dp+oh3xlZ8Al3ztjgg16xIa9mdRqjJ
2pdwe4UDUuYwJtpGbeLrvA4jCcRhdOIfcTaTaCBsQz9CpS4qq89zg8amjtuJLrbbCGYjw8H7zNcy
lfKguAVYF3SdkP/JCvA8Fcs6C/Y2zhOKRkNoHTPs2VrCIZTx2miBn5JRq8XPo3vY4iGSD83NbNkp
wU3UeoHHF2HAi9DMnxP9LAP2aC1DtsB+NxRnRc16Mfx25OyUGD98RDc9hLURxErAVffR7GqkxVfb
HSbblo97tyUCa5B46soiMFxeNfoqs1ZT9lX7yE9aW5MFIgtXKjtLgwlJLvOV0i5jXQTd8qq++Wc0
sE3RgxMa/PkiDtzTNkyCaILQvkhvM6XOY37RhmH+J3mqPkLmQemwWM4zxjK0q9f8RWz4LwMFnBXB
bLWBk0JTcfFGB0GnSGpdAFtja8jBIc1J72TI3R84X1nvzK7b3tUfCR6+FFxdGGYxduxMW5+ZOvDV
qUiGbTfJ2kyob9dGtZ5aRL+KMzWR8TMUhWJYoNH9BxP+waXmB2XkNgUtXky94KxGQ2o95uscuiNV
44o9UfrgQsL2l2ZnBgKGWxZ1PPLkr1fYfciRnls6DHUyVtGjHyV569i/1k09GNxPDaCp/IwQiCuu
OmwsYl/Ij8ddc+2oMAlNkk2yTMWjZUSaF23o/zhfoZxNy0VziomWqNS7vxO8fe1Z8FSgPK8Gggzn
bqEfvXgl0ZePYOwq2lsF6FBa2THX6BDqRmqCOGykNYgLkoYpmhNEHo/doWXhzQ2smTRhybyTyCNL
8EH1vpz7ceY9+8I7YQ93aOvgz4fTOasJQRh5FBlKEq+3TOBBUnHQlsa+qwxyCGsdfXpi3hD3EEzO
73CTBXWFhmp394AeMnYBjSNGSugDPsgflu5hSIPZVdavTUVN04CLs0FcjckaH5vK/i7qYr3E8IA3
ZKwWH/YfrjJjUABH+FSF4fvafdjjbu3ZIR6P4txDuSwTTyRpgAwMgYFqbZabrb9eE510Jl9i6EsG
h633WGNCxnaSWF0wuhHL1PUMHPkjTwAdWwfmyLAHDWK5ShTYzeldbxoTlse6ea135rkyeNgQxsaS
++TNac/eKcnJjcB12PaqeQ1LXUMw7VfghliADhQ3lBu4o+N3sSXhFmUAGL/ABqEkGSbWUXechSdJ
gIOhH6nyxB52dLqNOHsyav+SP9ru51PViThbNJUEQJ/LX5Zl817qp0U4IhbQWH0JFFEDI+0td8Z/
ZGB/Xj0hfv6eFv/zkoIN8hemiTHsQpDr3NoxqFqQBEjDDLCug2bGG87QokPb/7PvnZDbMtUWbNp9
UejDHPmUGdcPlQB0SeKbDUiCNk2u8S6y2yjUmzx6citfC183mjXqS4jZzxcCXbSeMBx9i4Zl9skd
08bcb/2j+FI3M2Am5VoXIImNSFSN0I4et8yvzBtnQxfUa6VjSDHLOfXPHEWeQEz8ylma7Tsv3qGW
/A/opfG+vMpr7bY42wwX6lPyPitAfpC6SkuJkPgXozK/hwIlNRXatn26Bm3Vkn6XoRPlzlw3GLd3
k9BRkDmt6icFYsSGdkD/krSf0QnVLwV1iS2jfXskyx5slpEqQPvTVPMQzk9VHDfxAEWHCGjKCFE+
IPxl2/lu0Zsrq5FLQA6nA5zalaNckBIb4euHU40ZijaCSEvmDa0zjUEDjiuFvDCeS6lSEffs9MMS
2Wwb1Kl6z87JYIRIMuyLcmUXEKAeZMC9bJa3PGs8M+u4j1yZByxLiyQurPaoT3n11rY13v8dGQY3
qDB9qkIgPyaugA1Loe3DDSu6EfEoCWA9SaXadKWmecn7yp82fJNYREcD2jTcAYVM8W+A4g2nsgSy
pK8BL3KbIdvJXJT0gEcB9FX6ykjDPPqYrkVdIVzI44SDN4Ze1pJew24lX8DdTovXGHEJcWTEL1Vk
XlKU/2TM/UphMG14EorzoFc7FGWIWUpS8BEtIqEaxxxsFcJYzCUr5UJRx9fbCYHOPvQm9G/x7BlD
Hr5NyrD93XlGh8EcyMkVAZt2kSQih348Jgs1hSw+H4fLiF4VR4WOwqF3zxin57Kz9OIkY6gkq4QG
PtVxAHvmQ2c4XkSCYal4AnI3W1vL4u3oUs5wb8+F8WboCiGcZQMfcuwkm20WJkNHD+K8KMzrzas3
AlOpg0rrYUrBEpZnns7h9oYbuJCAvrT/mV8J+d0S/tnxQZ07Jrn1AZXHROKLEmva1QlCkHbc0F+y
dV/piz8c3RisM0q7/ZUGzj/krt+vVsifG1y1Jgu0HZbTogFzrh2tKDWi06f44AdEzskVzSKk8h/0
Mk8sFCb/MtVI7ND3xKuyp9x1CgybDeatpsn1+JvnKzugHAs7aVACSuj4P5UQgVqQPvjMidSfFL9l
B6TVv3/uauOS3zxfe43jYeCwbkrN3YEwbxamHmBHnesmoqYQvFnCL1OeZkAbl/YamCZekARXrnEj
vVeNZ7cfwkbsnt8WM+tPIYAX+uIJyBvXEjZLKS7Og1l6lMstRDrg2m+xuvLJCQsjYQ/kQnvfT+jQ
dgU8CnMrzCsNB2IgP7KlJI1pTNqPipsr1WeMlIplOfHUrvxYgas6WOzeFenx/Otbvs/Brs0S8t8D
ehLRVNfWH9ha0BqynWDsUk5k6cEZRFdtJd24c8Znyg/1Id6mOzKH6zC5SrZ5N15S8zEHbUTWOCNf
3pKLOsl/lqY509OUjOz0XPDnOEGH/1Sn/VssbIcBJPHJwObvQytopPVX+jO6MwR2wLTtBgl9Pfmo
Fs4cSXozU2vvqO5bTQHeh5WSV8DC6DAxHQZalhPwmef2+pJtmSlfdtxNqN8DzrFFMCiSONXLCP0/
a+O6iH4PXGdEIEoDdj32qlvuUwjS7UHy9buiSu2PaPPOuyf14eKISbn7tWDSoTyi+sGjccowirCN
k0rZZ4fIsruKkgNJFHc+VDLkdJB4TaCV1A9rCzuQ7+tV3EzNxI/ZeP25UOEDjOD1ahgHXJiklNCp
B26QfHyvUOvhPlTPU2n4jVTtHW1XlrXdhwv7jIvRi4jkqpFw3Se4MhHBt0AVlSkzWb0Iy41/YlLq
xSRwrQxr6KLUocsQlC6vBKxaPb/rLWmTgsTxvOEr1EHqmLR4xVuUGzjVPGd7FWpi/o3dByk3fK+D
okhX6xBqPyVcDbLaMbAL0tmjGTDbBpREMZ2HIJJyo/Y5SeL1cHmxps7aqaXncMfzCPMMY7JlXrjk
oE02z40aw1nDPnRKQ3or6PJoVEl13ynzhfBQfxLax0FmsrwrJATDUKILd5e0ovt5deE0Tab/eYTL
sTLH39t74BbOCaoDD84c/jh/1qPQzxyVxffYQTcTKfUTN6Pwc/W7s6fk/ZDhAZhQJaZzaTvgHKkZ
ZYeGlye/itTCnb/qsI1iyl4c/sdM6T9J9Pa2F853u5iZqq+XKLSCeS7xYX7/80w3tsAVqMU7LZjq
hV+10GO2An4PD3MsqOu4Bik6re+EoqFE2tpDeKi/OysvAr3qsAO1xzDpuxMRjgEezK2ay6AHD1u/
q7jG2JiEV0QxmRfC2cOt2D9IfUy/RFXmJlg7XewaDiXwghLXhlTvvPm/86Qisv7wrH+u4fIydjsv
fm3qpw21M66/uPmDzCIlLRGj56Di2snfJfMy8T0boSIf6Kmhb8GD0Hr+6skdQG3MHdLSJX1l2HeB
IQ7Z99e8Lpj+cdRgBM0j1z1R0H3wcKLx5OXu3e/3X8W9AC00k/46epcYT3GLfDNSB6PI0FONEPqT
14UyOrxRKvtp30I426yfCzFCQviTw+8LusO2a6/Dv7/TOfMSUoQkoYWYi6GwXoetGHb2Q0+nKSBF
i+OO7Zpw+DOeUOVuv5wNc7HAmN9kASL+nw8Q/RkYI2J1Fxb7v+kiLw2i2SRjuTu7kvbOgRI6ItI+
dJuFpj2gqN65UTm7HRLQkk94qdA3AXUBsSbRoWY0iC0cWaHd6sFaA7v9lP+53cukJXGQyAj9EJxt
zTOHqkXQsMrxSaeoShVxJyQ2VqqRe9x/5VW94VsdhifIszTyudUKEjXCq4wyspooDGwaqEHcrpya
cOdLA6Xq0sVL8xlAfv6gCjNcgl9eizDkP5LzofaY2Da9xK/MI/rkJB4uMNT94KP2nujLe9aduB8G
QL7er0Zn9OPHfguC+yL9l2lp8LWnJcfCk6cw8OpsFy8bbHuuoYA+gE3zK3zx9ckc2/qOY3jmhnId
EfRJSMXuYk3OdWekg0naZ+MSuvr9mBCsrg+OpZqcldEcI4hhVC1u6nF7bi42hgTh3qC4zpxmB4ca
GwIp0vZrFF6Umb2FYq8W/9phFentP1p16V2a/Chp2v2foc6WvL+Hj9lgfWMVp9ti3zr1PkB4dnuq
wfqb0Az7co4/xneHo0mB/NPw9WbFlbU91WSXZYuB//Y7b/wTVSonlYEIETXMfrI3BLg+He6do6Xn
1mvYTmR9dpldSCOMoUdM8G6nWDUH07Bw/cuxwQwf03h6uRa2Hwx4TVPolV1LX17V9Uj1m0d3zm1q
Upqn32f7yHxRxh0sH+wo109x6m5KwjuZzAN486nLr9+nkgEHtPnqGVSjlQgz2hZcEczuiX63nRhR
z0u+YK+F9JcOp8vD7q6/RfSnlxjsd9SrjwPZYlGaA6DacSSqzs604MRsoShAWv6KF/td5m2wUiwp
5x+eXrl0SYi99i70gcRGx9M/IaMDmmDK8ltZ4w4YfAJhAN7bVpwj2/KQ3HKoYCzLZtQ0gzrm3MLd
YcdQ511cUk8YyUyqOmo4exEjTZLEHAuDy6n+bckRhU2x6qLhiJRkQgDNAxc4+qgr9JiMKY1haV3d
z98yJ0AbTXb603BxsnC+A9AokQ8iFeUYqZl42u6DoVQEa0MAVRLdTINSzfWBqV8rfMreSP7rMs9B
fiuXRCBPErNbI73Lw6N88ZS2QbZBiEQw68AYGpYbsCVuftjq9TslHG0L7qo4EYHVZREGUPLstFOW
+QPHDnG4J7iET5zqqBlzcM3gjtuz4R22w24bUMiFdeCDdKOpTkcvd+N+R7rIHKsn2EnE225p5T15
tsAXd+I+It8n8YccEEOhaTQnc4TWAQObuiwVIeKWG7C4oxofVt1D9JxCxjEDsya0h9CeHgmhoLsx
Aokxao1KmIxUc8v8W4U5lQdx4zjXRqbTjnj050ZgVHrrMkgv5IKKgtjpM+6LXihQklA3G4/vaYrJ
Fzx1bNAILzmE2Sj0ofFIvaNOzI8rWvYNmple4cEo4S/+yceoMQPE7VNC8nCgH4OXD7dSfRuZdLMr
7fZFge3N6tltH7CscRNV/PyUBlkpuBqrXmlYvHhZEBym1acITRSAF+nPLOnkdzu8p1c52J1WiU+D
Fn4FYCVHuZN9UtmIIQIf3Qd9GF0eZeMP1UFyGZ9m/JsfpY7uSND1uphEeD6o0N/JN9urCQh8QB1M
xzdMis8gS8EfN6BM47GaUUiqyKDbOp1ydASn1BKzjoXc+J5sKTPsffjQ3EIOo9E/eP0FX7G6XPYS
qgrzWEZNZuYNbQsO5FAQsJtzVrgWOi6KVVsb8uNVFXoCpyS62Qd+bMI3g2DhXCT+/RXOx88qmgLB
Eae2TQmW83wod35/Y0VGesFkXBkLxP22kHfrKmmRMdpxWZGpXyuuWrv5ImKXrxzukLdGs+qU9NUj
5kDZksyrI7BPsrhydOozItz9DCtfVbZj7Ig5I+v2HFKFd5zDt1wOhXF2JMDkUrCD9l06gTTaptt5
bM2cDs0vy7DTBnnaBg9n1GJIrGUzW5hrupmlYs+8XKGXxoSP0R7oP7A5YBBgtXVt4uNgz/8ieKD+
He1LS++GNL1IwSXCsVvqaMU9XlNWiisSEG7PU7ZcxjvF/gSXYJ90spljTwvF8iH3TWbMkzM425m2
+ysndAeBD3H307mmIEGmmbkqYA4LHbuwfBQb/ep42CoRcHMpxQF3mHRHmATJXr4G5EHfKpQYJsdE
g6bEUf4uVoaS1nF7jOtu6A+QOFDI4btF0Y2ipov771aY8A+3Um/tj0cgCdXaK6AqFs0WtrMxxEZK
TBk6qOmQV6BETUYD6CEViAEsFJaVOWlpMhvPzmGKH38ft0kJG0kvaDNzZ62yO5KpeX4kjeF4sM4n
C5BcD0RYck49LTei34nLGMT1ixaR7vJ969oW6NSYD/KidW4rQXPprT9vGui5bTIzDRHVRof/V0UZ
1irxh7tKFnkjNhxSWKcTHY2W6VUFbKFoCwND+z/dgnsVZ7WB9s2OTvYGTS05hibPWxgajm+eFs5k
N7uzQIgyLGEsTYclDYy2ANRV7nfERkIURP7g4KWit2bfFp8+HIjwZAaKeUM+qE49klwXvgJganR2
svdPKKac5F7jmOE4Jcsz4DcsRi+V0u2BREiukLgJ9koCnuh4kS+T8rOHDkm33i3707wULxfR9ziR
tvVmHBY4I2uPzxm3TOT3ZcVnaa1WdMuxDxzqcArWircjy7fhMPtd/YRsAH2El7ATisqKzILexFxr
Vrn7S/SvlMYzJ+TQ8a5WoFdOLYBp7Dxbi8LTFFjtTgGzJysfhHmQPF4Fx1GNXR22JF1VPsffikhR
z0kJJPPe7O9R07qU1cdWZJLk4xvb+evGuwRrjWTLVAukJJ9MlSVAvpEP0B471DNq7+AyyAjeMEJv
9RDJ7QJaTNUveurDpweooMmrqukkFmCNTOLQL5CpNcDB3m5dj7s5nFJ7O6deHTmxYYBaMSY2tgDr
nHMKpuUOyq9UVm3qMIX8Ahx/7mUgBB1j22lGOpYzL9fkoMVH0qkwkZozag3pDv85/gk/BhsMwbKS
ckml7Cv8JoIg2/VNrAjEyM8fSyF+x2i+NdbuaXcVdGkm82gyrsSf3JWwt+vchHKNDm284RET9jrQ
OhjhKh2Y8/3XcVcUvbwmUQJ0mrsNUeYg2anzqntB6h6SWHqMgvkVdbYr7b+bzKBd/RcNRP94z84z
n2FVH/FuRpIRYe8Q+8pJWQOhBg9Ppkk6+rGmskPCi4LPfqnAhTSnuW4uMGl3nkHdKESkAZUlZplt
2pxrOnVABklKXG2ALgLWpS5jsoPzK6tqzHRrHv5K3Ecm7h2kS81ha5zQKppubtD3peb7nWEbcYG1
HCOmSMQ76DQ77LfEhYmiLIy07MPlAz2knDnymX/MyN658d4l2uKBPoSzpuZbFWy9Ko+Hfk6RUzec
6FzZQV123s1QCVmow9lqO2eHnL0PqT+FQcbRgkW0O+E9Kfxp7gFMrTkTnLTE8vEtbR7SGZ94v8Tc
GSqkm7cRBjQmE+atKe1UovnX9whYS9B3YOfahAwtVzbWHZg/kUOoQDRkgKyOqhZAFl/h6hKJLxXF
IDRcjC6HHvskcpD41BvcJF83Ngm/XIle5ywCPMzaFk0QrreThF+AcW9cS97dRs9sJopySED/qypR
m0puJD8Mk1b8ALx7Csr9ZG5AjIltcPuBapFXKg8I7gxXHLUaB++KbV51rYiQKMJiROZ/PMMmHtnZ
/mTkNpVR52JiQTRcaIlzobh9WHl2FHn0fs9RnrkPD/GzQnBLhtyZh7zQbm6cVffzt8R6EXIJ4Sw8
YAsNcLrM938TqpSfMI5m989WUOql6a2HUfTwOIYTiFmV2sR31AJhAB8I2+ul1aAmDl3sZMRdXVjv
uCGXeS8TG1bqyt8DHKLGSmCxecAypl6+upJnZpFkZJbH+bjHXhdUucwFuoh3u/Tv4Z2L2dok0pXi
a1EJTEVBCvCu3A42w1XDjgY/P64drHvkm6iNId+1foMAhxc9XeIwSdzsoghZXHMDUwPZeo4IKrz0
suUlYaOLbGDbvjfoSJUlz96C0aUx2ME8v+5SNEkNqDfZBG1fjH4wqUo/vx4wyqVHz9+N00wu6ubC
1wHInCHxHL8fZHQ1FIBJy4NkNzMGNRdPn8WyCNyVqANw1+L5UxaLOy4sqK+UrOLqBpEtfLm1nha7
3SPbjgIp2VIVQd4sHDpWqNeNH1bpcKMvhcmv9sp/a5Q+uJlkO1t0GRSpQCsm0kty4oWSe7UWOQYH
3aYQ8HqD/9G6Guq64JaQJQwClEVfeO1t8X6I6RQEKeX5xyuE6gzC8p+TEzMgiYNxgSPwK1BnKLhX
5KVDe/aU60tPD4PiIR1xY64IcZAs2zZu+obupAukdqEWBk7vbNNOZCdqDf5Pyk7CwL97P/8SerW2
ptJsS0f6b9MOlv65f6P37OsHH833Fgivi6Iay+GPM/pSlBtlbMtVbzptYZBuuf8023R8/L9S/wJB
uiXdR0Y4wBTK9QN8cv/OvZGqBokUknE6QMadR9iAsChjchXEyVrun+5szNYbyHgfXkzY+0Yg3whU
9gBm6hcMyxJI31u1MnKgat9SZhV1L2Lz4/n441DgkQEuP4GHW3F3dnmctRXUI1cxuPGWs0qKs0u7
GHNjHk0ghFH3+JAsaLVV0ndf3qc0yuXZWKrHlkdd/k0k8BW2S5kcljEhqKEVzrwZ9x0xDbQ+o5RH
wZMWgH7ZJBVUazVPipaWChjAWELZoDxMO2InO+XJNyC7e4siSlunCvSVLHBzxiCjkPDCcqMr4KWC
XE+oVPGCYZxODaUpPdgvMobme91AsG5kf64A+qwzQxiHYl87qqVWy7BC0hJNkV5bETPdCvDjaMlu
Rhw8PfuaDLz/OXvKQ8YYOyBslrPjNDwYutN7lk9TJVRizndf3l/iQQTUeyQ+c5HKXYTXuqbMKGUH
Okox8rN4wxcGHqVN8dmKnqNiw/CBZihFJL9K+xzc7cmm+qDWGC7VYYGylyIMHzV57C0YfOcEXZFF
GHBvk/u2blgfTFEcVt9gFNJKsyPNvW1KwRz2SPYXzUFg8P35XWggSZSlgZNZERN1wyppSN3O23ef
CiJu57gjac7sAFqS1m6BZF5iN+gEcegJJDtJX0As9Je9IcdKNi/Nw1XTQs8hqVw7FB0MoElbz674
LSdFYYLco6PBGE8VhV6LuBOb37Agy0qkncNXGXA56xUBIhqWRHrcywXbYzRb3UawP+3vESV6V59A
W2NLR9yV/IfVRYVBkrZBK0dlCz4WSRohZecg+4r8NNKD1gfuwPYql5b+opdg3UXD7n99L+ZTL6b4
Hc/fd2VfQpoVWr9xpJwwFepDgN3HucTS7p+YLauj1gUi1GoGa3jZzFJ66T0sVABCnpRe2gKK93Y0
p1dNjJkzbyCXI1L22kltmIwuV6OvUt7HptOe0E1u+FgatsvJK+jnSokLyDT8TSTjSxBz6PNO6mt1
z0KIMmkMqgOpzx6e0Cypq5ISVXBzqgN52gbfUdDcRDN/GkLS8Ogu76WMJn0BPEFa+YXzSXP+PeiA
Avn7VUnucLYENZOfplGvENE8Zez1Sa0REaIAf8YIswMz+P8wz6uCraVR1rSMqwYbL456BPTzwz5l
XH0SKlQmBo8+Fgkwt4Xc/HbfpbFHKToETvYFQwKpZP1leE5VBwcaobvjwOmo1/V5DYxL7nBNnnjh
1SHsfJFLJRLGUVAFeP26otZk/T2RbFza4ZRBnA9uDqk5qPotReW9Ip07P6vzYt9bvUloxZSmaFq2
ILoBu4klbQtyc4tF2T8xvckZPe8NIDZcr0GmHcI3FSdKyVB+Iw6hG41Dys7v8Fl2wXcMcZD9/Cjq
ZRDu2z6tgRw68+8xwt0PQwHXUe6Mp4l/dAyArSEqk3Tp4kIUK/6CGO5TkGrt7BLxluHolY/jyC2w
28rOOyjJJHJ1R2dkrs/1TZmjKRTjd3iRniHxV8eaf+Oe9FcKVIAIINeHAlG81R5ab7f7ijTvOFRQ
+wdOVShtepecxHYNx/CIdtAgiTFfjEhj6hX62o0MbenakNWKpNFgtDSnOtdkVi0NHpqLLFfrGoIO
uGUaf/rEfNY6VWPCVQzVRs1rf2fUZjVr7ajB6VvLk7g8usygP+cPjyUnGLSgR54+0rUdynM2Yr4w
02JKqJYO5YXBlwu9bZpg/WHSaxJjn5QtvNFkIf9ajsjyMCIkXN1ipIILlhk7SE2GX9yhxjjRhi2I
5oRZ7EBu2jVlNyQpLPT6k9/w658w9VkvpHulLnkuTemdtjRXpRYBUBO9JW3sGZa76zmQjIDy9hkd
d3JmDbYyJ5+ecpbM0G5rbu6BD8TcYaSrTT364h4lepOjm2/J6MGVvXVTEDROG4WX1tlXVmAOIpfK
FSUR/6wiW/VFPBNqaT2RbwxDf+llp1VvxFvudnEL8d9i80BrXJouP0r/qjphzd+zRD6c0MTXUypu
O5MVzmWza8yEFJblzGtZAc+Xj0ejdEiDSKSmdgKxkNi/Lm5ljWV/mv7Y+CTaLd+peEAzyLhKAx1+
kLzX0RXZyRBR7IReZIFBX2fpYVki3RB9vbqtFbLnP1uIyu//4P05iL0p6h5+TKkxpE8mmd2Lr5WN
AQtbpP1Vp8f1Zv4dLIBIOBLNcsrUHyaDiR5AwDq98XRUlIazvD3feiYieAH0KpEUYlUS/kSAag7m
YmyACELLyaYZbCZnHzQ4k9PVB/EXCdR8PPX2oTsWAmLeleRe3r/fHaYVKlTncZeDjsueamiTX5Nm
Htw3WVwiLkj9j8CyRIgUefNPxE8I06HDKLWJWQkVsAYJV17cHHJUuwSi0W/rg+F/HaxD6CZlP5qs
h8Jx5uvqsUuaQ1cZbEeFrxVqktxkLQp0gs1/Inj6ORt7361ckKI5y5Tb272v4p76sAfwOeNPfJxq
pAI80AkMqJ5hKVFzF5Bi1m3TXx5xy8jGf/g8n317ucJPr9R/gphNldrUdYWk1d1wYlRh2aRCE/xT
5ydAQ3ZR7BW7Bg2G/ViAO5v/SJG77lg9j+nxCoa9xrKy5HQLbXVWQziaB1F/ei+wBIG/McHg3eoO
RW8N93UyI7OmSY2DcAoL52Bcq3mnq9zBSHOO+XWVwAIngNSt4RdxJ9BnsMac4VLRNaVYSoh1MzqN
6HLpXVJtu6whEqJeDJlX3XXsEWRF3eobr6cHeC3hmSlJtzAFL+WSlKvKXw3FAtqyDohda/KTFOqv
/DQeT5CholcTYokfoGBFubu4dkJNn10I1FOWvByqtMBdhF9qNqR5A+dP+tNSl5e3jOe3Udomk0Ax
gNjxsZ7Z4ZMR3eJje6hVQ+wNZj1lPgukLX9nFGgowTeVT/2eagAcWivLKf2jipwMDaCxdqD1kSn/
9WLkZtLY2GnT4gUdJO6EweUub0rkcUFpdkdTbfZ68hhZGpdFPKm4JzW0qa5LErKO5MWCPyiNg2v3
GDC+hn93T2vzb05JtkDk9uOze4+73pRBhTSX7hbt0buJax1CegtIwHJlMsgcwgGSTLL258t5x/4j
LtVYLj96IO4mHLf0Dh2ZyzIUarI40rOp00VFCE7ycKjIe+WilsjPWTUjxwBO/l89ij+R1QCKpGPH
GUsxVuEwvfgZiaUQgCITzKPsTbMPmCjlBJLfyOPOMHbyq1XwPMXy7sxG4M7HTXfjARXtkWDarcPg
EvGNEdp461fZufrL8YnLJgQU8MtzaXjfCte0cuqtvRUoHHYmuEjg0xYfxjg7cXwoAFI1hrHC0S5W
Q7Oa22XQVf7dSJcUNJhe16KViYdldcXWgfjILybh77n7BmazCLS62YN1xRYn+C22UpUP2YrE00pW
/ywGdFedj4CQHE1IeS+N9cx9aqTpzMXaOoEmJgYh/jGdSNqSIxpAxXTsGPyDx3xYytHUQ9IANRsc
yorwWdvK4RmdYmwCSzVWW7hU1ca/0GaK/PZPOJIyK/JHF+YlBQHKSJQzQM8mx0UWWHn2d5m7Etvc
amCC86Hz3PYj88QNISxMCeehk3DlX+11rngl3uNmB04NB4T4CaMOEuOydQwpdVa4L+2rUYM7qKpj
rteWctopuu2zljbiu4U6MEtKTWRwvdnXSkRJQOGDCnI4pLi1UaciVegPhi/WbsswC8tAT2zH5xQT
rZpcqlI6bHW3kgd/7BW3f0T3oaWr0QIua5ERRY+lR8PiGN8C33/hRxssCtg13jApqgXT75Pmk4AO
BBEHLBWQZOVQZ9ctnBuz4yZ9/82wNIODnrJ0T20MuX0Is8o/x0Ng/CkFNkejtZSJyhmHed1wMsM1
aUqkLSIuCU2jh6FdLM3S3u+J5uYgnizlhZtQ75Srlqa7qh778HWETRJkCisJaKtCOaYZLNNic7Xz
rAI1E+JORCFB5G88xlFm4MVYR92XeWAiBxofukQlrtpp92bpEWWBZRQpwO7gTtAfgMYU9syXD0/V
Y6KcZf5i4VrxVAWWHaoYrmTNY0ZZitOiLWKcGtDbpvTbeV5R2O4zkwGZsVdKlp0h6MIPpmVHiHHk
i1bWjfPhtsSwG371EVzDV92u2GYiB3If1scbKhARNc32mSda2QeKfOZ/2XQIEjXQ8ZvLyBH4NvyL
mWcsOeHcGNZkAQKHoPV5FFSxqo9eLNvbXcj5/1oguO75TTEh8J3nJyEM1uvrdDcecFMaGMS/9naY
uub4h8+SsAuQcYtg/NE6qsTic6q+hPfKtEvlFub7xfCj+wN0AQR0XL0Z9wZDf1bhZypLOAUocDMV
Aw+zBygNR/oM6LNmz2QDRwtd6dt3fpZw7zp4OukQoM6Wozhg0BTxFUcPdidUVkSKPOkmGvJbOnao
OVGD3YK2274s94tQ7psk27FiwYZvjzLOH4KkVqwfcJ9u23G4SL2sTL4LUXi4k/voZk/dcgvoWgn1
MqAtaT9lVYYY6/daoJE1iQ13Jd0XQnnT+xAzfVsZCm6F8NzU8ZaN6I5j8MKwbiYkrI7QWZXHoTyH
HKfnXbQmOEJ8kMCC5huhSD10nd0qrfvuRKVdirrOyZcCqiODSQ2laab0Ntty+ArTSBrxcVdtWvbN
zug0M2BD0m2X6qN08BoYa2BRkgrFPHcJd+zbBVYurdVKieV3gSj7cSbrd7aUOJuSsMkuZX0M1AqI
4379u8kjQnnJk3irbfJe81CbM+eMNkaeHiYWGkTvxTmWlop+awwu8BXWEwRvIRcTLTvxsrl+3JTM
6wCj9lTwDUUx/nrpsvHiJtpUx9WDL9PffDWbEXPq0GOFW7UBIq8d1dtl4BoKYNUWka7Yjo4AVbi8
6cmAuNzTTC3u4Zw+8BVRZbxMm8MFl2dmo8d2J/Vc/QAtqopefmwdu9lgvW05b0VIfS8KrVkOfiH3
8+6Uq6h4If4IoGVSiFyGJ2o48EdO03F3OWE8IZHmGcAkuOX6McmNiFzMEU59Kzg09DuHe6n9eEAn
T/f4QO/AGdRxWxaSRu9wvR/AynVNWzE4CbchhGVRW7V3xudMhlptJEaHb2IZocHDNLTerClV2MZv
uMxFX8DPfCbayl1DG0JwhM4FNixe9ksnq3h4O9ziR/0booWc/GxeAeRMGkEzkuzcgxDh1Q5y2K2o
Pd43bG/kxjoQb+jOnrBsk/OxJ6bMSmIgfQmLf0EGS3qKgfQBJiHxlTJpice0Fyshp7Uj5qMZE0Q6
5zn/rb9UlBar2019bBxguN5qVb6/0oyM/kbRomSt20BvcQfkOqr4tNB/bybRffAfpVRJfZqmYLqV
Iya1MnkCFUjbYdaO/we9pGi9KyrTpiyVUt2beyzC+2K7FE1cXAUybeUB9rsMLDNZI2pxblBzotzO
1TUAn0yXTwcBLQfWtKhl6+ekJh6A8twXWnnYA6jYYrQ+dEcN93Y5iwYcV+FDEPBmugvQa/sDache
1tOraYPzPu2bZ1p21qhs5gbd58Sf5vqQIMiC8T5bdvO6YG22xZ6Cv0GEKOvo/WhCQNKsx61KDfuD
HvmIfDfm7TJJaseUJ0o9/4uAzevot+dV81s5trFJWJvFHepU2IXLEvwAkLklRQVwWy9mTSVnnUT1
cok3aL1ykw4wAl0VC8dhh0us2HwMcztvbul5L7Dku37D+OHZFmaBOLLg+aaFFWm1H7D+9dSFsBpk
AgCzqQMF4r0WWhrPVoUX43nZcUSxx5BrBY6q2BjCvhZlP96MQx2jyYotW+eC9AqtVoKjRekUw67i
DL5lmnKNMuuaXZ6FJHGp8qD6GbaTdI+EG9RfvPKQsG8tyvIvYAUx5Lt452pbVOM4ss59F9EdLLjy
QVJQVeybLvLGFeEGeHg/yTYhNXtVo7mx2mzgyf1awdwVbHRzw5lDl96JP4Xf3Gy5yuDIKZxJcXRN
wFOtqlgg1o3GHiPcG99hZJcQlp115B78NcMZu04AqZdhm92pnSJfCmcvC9qLcwlFaTlKbFF4TeLE
X8P//buX3pzfk3+jmzyUo7/oer5d6xZ+m4NABIAOGXAWH9G+XYgs2tokMcZ3F665nk9h6YPAdmPM
mfsvr0UHqa6ZKMT3UlSdo25HPQovT04Dhqi7o83vi6DwQCbfR4k4Sr/K35RLne5mF6XMXFOTHKTL
LkNsYWS+EGsWd56vjeDJKShmyi7KroQbxxZmVlsszLAed1OZcgMSBMAqgWZm8C4wnuSCCF7s/klU
KyguupN/oslS0AlPuT1DlcNeZRzw4jYBKZsnZzHg42WuyP0NelxvfNQNbN6VwIGZKKU/CAEEq9Tc
pQ+6AQof8YI6aZRFC0cOuK8K20s2u5nh1XNqXWxyortt9aDp9cMJF7v6buFY+izUgIaxEXK5vSJB
PEy91zQhpvhVtIjTk+45tyKkY89k/sF8vncnO58Xcz7cK73hvjA+RBUM0EADWtUnIoQ9nQOZCQ11
Hz7e7F6c8oTgmpp3Si9hDmP5ZckZPCLjf/ePHD6s0dwqitFdrwphn50K6LLTzxyNTUzVUNkAiArH
mJ8y+yfcfP15LakoM+EbYd2ek7sDpDCYSaZVlouCmU8KYrnS1WczmN9aw27RuiiZJ0kHXEmWeoLG
V8n2GzFPTgx5+xBjmU9HEEnW+w0NillQKbDv7eK98/Zx5FoU0S+NuHmpbunWEzMiQ9hrlmn/TFza
4pO408XiAu56qFU6Hag1VXc59kTqZRe2rI5hmr4kVEb/pf7LWfMndW541jm1tsKJNILjJZpGb86B
LrFUO4qAON/hFFQCQbMZf1ye44J5+4eqKdZLViL+464ud4+2w49SVYSwYkh/QQn36+kB1xmr/x8s
s39y82uQMpRerDcsyuq4sHDXo4+DYMJzT5yXcH2gUJ/inhKxwdE8f9+yeq8b/vTWENN3ldvasCqo
+JsQLflcnc8AAZn9RZBpEikhOtRNS2qVQj+EUbbIRGoy4JiImyIHVvey7KrIhn3fTTneBCa7h5jQ
eUhsZFf1u2jdZSahiYt7tbSQ1NMgBQxR7SvYF9dC8cIJ353v6SBG7RyYxJBWCsCQGXLuKlCjkdGS
3mfn2ev/tSt08y8o5J18xymWue5ugHyJHdhhz6ItPDr2RN30o5m2tlsD6aRYOyimFIsxiAT574ls
RcrJ28rd1U0s1G8eNsu/3BAEGAo9LVd7g7IwpjP0khi4GYjhrYKtsSJlvR5hYBKRRkCvE++RVtmA
lyLS/oqObUO3vPOp4Dqw35nTle1mnmKlZ8MQTQq6LR5HKR8Txj4+ATAwVYnWrEdvsn6LJgPJGUF/
DfHxGB2Q7aorsaCSf8yegViJjs85kqBc3M0kK+9MlGDKVkado3eCg61w2qX4V2V54WjRwis+Kqbb
XZQReqzyJ06//l2074Opzyhsmk1OjkuwRZTqgizmOtK0GoXOXDA6g8vGtONp+mDkdErcT6azjx1+
QIeORH7s2VbS4QCx4PtpFIGWK6E1T7TAPD5TWARwJqJsV5hIZvUjc7UNMW6lakT4tqcUioiOSgWR
DfH51NIgR20R2N5q692a9njSocxxmgmqLmTOYke5FpeFztgTygrAqKJHCyb2SZRs546nCcX3KJOI
kPmkDn4HtTjlKxIYIo+tf77zQufIJ33zvwZVhuIBLt4z3YVtbblAYzmyxZEKJLYNB7+5/7Z/otOp
DUgL+bNYghmqfFY8KeDpn/kx3f4XVUQeHgIL7/nvBRRtOx/HDLGEEVaLZbyNhXiek+TNebe198o7
5cTCe0UcsG/0LGDqb5XHxyDPHDjQJ8Rz5v13m3ChjCnswdBkReN2mUxce2hqWD0C4nxcJX9Jf76U
ZJxx0oos2KeDnotWayK686Pt991EXU4n4v1At02IrsTChTTibjNvLpbNL3ki2JL6TRoUyJQSapUO
rOxMYaG4LbFqXVIkT5dhmmyRFTv6DcKtsglht5MIjnFrWSYi8mpmnaRKXAuAZkBSRhrolBpK5nVQ
jaovHwU9vJ7g86hpkJjV2rrlnabCI/DNAycYwwAGUxk7m8ZJeo72x3pdsAUiITOD41CFkC78k2d/
BLVdCqffeoc6s+5bwlVSDMbrI207Hifd9/hsj5LibEmpLx4F0rYu8+y5Ozv6mVaGVzFhf23YhOik
qedr4N8xDlNP2/bqBPiW/bvXpWbSnZaNb/qbfJY3Edgyug+Pltk0M4OKZ8ieh/QBA9C/vz1NHg0J
EXZFTlrr+y4gfyZkgs2Cob48zKPXNsgYl+DisZOmh+E8ZgHVPxDY1FNJAylO/V+Nb+rPNN2zoJBx
yCyCKVd9F6kmvoLHgwPW1CmLAShPfK+QU3A6RYfAjqJl23OR0b4VPMGcP2ieajDRv97RCfPb2xhc
dNJxr67zot7MUiHnunHtqTf4nUEUA9xlRGFhibFW+sXNFSDjn8Ohp1gfviF5Kdm5uOpDsxwijV61
VdycIrTCB7sduk2DlMIEzfMkf14oV9ErO8zZntMt623074UBB/T9At/+Crm10ZFFMS1A1HJurb/e
AqZuixy400Gr9pOlrS2HV1M0mAGXvwCZH3WoOzrUH1gWNkqWwJjxgQ9Z9+HSUbKZP7XoY98BIxUI
jbJJgyTx5Sp65gVf8PS2u1VGR/fBPNW4M1nF2O104D+K1o+pKJaWdJ6gqJh1WlZQZNkFo+RcZgqS
9yuSXtr9NsP30xGTGP3frHQXQR9Jk9wk8Ct9muZSigrPNeNxJ7giiZM/LQ/VAigY155HxyCINDBB
/KYP014qDiRegKb2lESzoHFoVP976JzgHg3dO6ZTyOG4+gQNBuImlGKxtHe0KLDofixFx1p1eeti
ZOavYaWsMdh1SkY/hh8ZkkhoaJzMt6wJQP683EKDonVlduvEZqLuXBY6yMVCwmH9k7acDsxhHf6R
aYz2N+xw77T9fMtipNBidFhCke+CufZewDOoOVHGmewK5h6ctGMvzHaYbucULeLr9Gb/LJSmDp7a
5K7AOfHUsuobbOCo3QNwek0KpteyWy21ktjmedbvOSi80WyMqTANxtZBZKDdcew8vOqteDtZMoig
WGdP+Y77AtW3uqKEaw4G6TNqKz4wRXVTiP7LxMua7SYz4ZLbugZ/CfbA7bFYSM2UCqu0AJTjcTO+
OXPgd+41UHX6ecGGtb2EZg/AT+M7w1CFh22yD+QBEW+tUCP6ciLk4pmU6ZtL8afQD5YM7syzb/Vw
xSGcREXErwV6r0+K2FpzznfzfByK611zgjh42uzJfbeiXgUvGaGaMkQJUDzaEJIF2Jd+9OFr413r
+fKm2O2yh51o97RG3Mgd38cxS20wQUtql27mbsDnOUNvZmCmeYJbsMRnRDe2M4d2quZ30qf1my+6
t2lKBbI3tGg+4pv0icP4LYaO7wkjeE3H0ZG9OcmZARB1nCWdVBHKRmhul6nMBM9g7TIo7a7AR0Zi
GLxIclEw11onT6YEmCBKHrQORM/nGYwN6M7lUYkHCbC+ksc+j7HgbdYP5mTOK5Mff9iUSo1bjoXq
c+XOd4C9n0FjyZF5a23PUjeePhpu3T3q0ReQ5J9mcQxppUaT/PIfmUQOeTMTB01u0PDLIdkAXds7
QgLPPm886cid2Gix8+iim05XMQ7K54BTkewFHw1iArq+pZYoS3dzQUcFxP5M36/0WRab22nECYxA
XtSbS2Egvwo5HMLYuBqtYDzNVuE6vMbpnpkLt26+9odQHb6vL+/K4wQr0SZPTUk/7YLDz8UWVlv7
36hBEnZd7tvRuijvGIX2O58OYX6BDqvfnbSBPwUk5NtGHwQ4L9yh9oZbVUHfO8ncYdhiCYBM9Nnw
FRV+JxeEcAxSq8/V7zi8LbGLTrEQMedcR6MnPpoDm6BLs4PL9vCSFFE0qlcu8rlhioNC6UxD3+Jj
ibB1i8k9LjMYjJrNZ2REdoemx6q6BMr1Ovx5k/UxWqOyNJGy7fu0t6rMlGKWbNfVBw8/V8jY1S56
4HfMK5DPBVDmLlI7QpNRc64zuvnk+yLHj/JxP/YlkFj1qkdD7+xN+6pcjLfO6Z0vGZyZKIHhKopz
Hxny50cet+WLrxeQCwRsDx2iBecKfiY8inoSro14WBUsmV2kVd98FmkY2LsUH6tjZzhtUtvUpEgu
Sl6r2frAvGuW26voRQOG0qCtPq7Myug/rxwngjhaGA54CNKNYU59wBdbSVulxj4PHBcw+w6QAF5O
aws9vccUTZrKHafwq77XZbuIlh2LdtkCpzufyR43GauFFRBllCC7XKveGaoUpaO3NfX+XmIeGzzi
Zk6Pei1KIzZ4hNUErNj00QvkyyIJQ9GQBHZXlZ2+YFVUFFTKW3rElKXUCPjDTZ/yxcHykB0YPlcY
s5c9YbwL0+F3noT/SBaWD0Fk9ccjqEyIR2psYrH1wdyFXzbnj9l59VwFCB5Mt8e4j55kBdxNAwdW
qKcbXALP9LP1cSDjJaV7G8kPSuIuVEvHTGag20l18QPNaruB69KdFdxkiU2SSEts12r8l+06NdN6
nypUcMZ7c+pmAU/TehC/S+58ydiSyMxArt/h5F+n5szmMEhoWx1FMTL8pxjNcqw2910F2qI866xS
kvOsz+RmoSgMd+34RqTfdbzNJL237lQ1jbRO5+59rC/9IkwLQY07pzU/AmfrHnnmwGL25LD6sOeW
L7PcRQTNTe8a3qrVjCb323fS3c9ymSz4+5sx3E0cNkhTGxI5+fGKy/2j3RQ0LskP+UB/WOieKRIV
P1O4N2cguFGhd8u1+iDACJOWv9jPKyqWx/XRzsUjUmHMZQAZsuBrCgfi2u/KzqIaVHwZtHv07tiJ
4qwgYeXlXQdt3S5PvHRLkKA3UuV5gqW9lWMkMgQhImkglRrlzCtiJOPzEAD06oKxFZzIocUqJHH+
LpHS0SMDsOxXqxHdGADCUCoTGsEUpXla8yjU2O8L76fJdNgXBrWXHwnm7AeacBEUGzHotqOxr4Op
/MKSz3OmpdZ1Z4MsdYLE44FFaemVRgjHrD5J4EJyVAJGnpc24LwOMb9+wixvUQqOncsakYbgaNUD
9zII2jlrPiqhfsRrAtVR5Bn7zqfYAFLrdCgqRoH6jihrkXJX6PKEXtraeUDjnmi+aoaiOaD5vPWk
13wo2ksfcQVQnTCCSXu7Xn8xeCDngkGLc13FtL6DgEqKKwy+dv3vuyrHo2jlnEWFva5bEZ+PthYj
/UY+EoLfvXcmFbOo2fcd0VslUgHZ49iDsv1T+FIfxuo+/c6BOmffn5qM9CR0BftHZ4ADPt5oPoAq
04wjlYVe+2I0Asfd6WJ3o3hNEi9i/9F4UA+Sklu8xa+7wLRlL8P2kK+1sW7hXS1BywmD48ry3XgP
RuFqmMs+EZ3IuwHrSg9PqMhQ7s7LPGHHbFoACmAvetdeaFrornHltKOFtOFYu8cA7wiZ716ZV6mn
uWgVpjuNEZyhGdXFjNO2azyz9IrIvcejTt7PRZqsSG/9kKrLDrNWh6MM9bsG56f2bFYaSFOM1Tcb
bCd8JEpUs1dco/1wou7P/+pPS6g+Q8+oIPnO+D7BQ3cFYyFb4FeycDhT2tdMLOGHBdKxWPLUW/Gs
2f/8iybPnOHZTGiv/UpTicoSOh7NWAXBjz4VaLBuyNWpM64qoV6WQgxdcTncH9Fzcnog3fZnX4mN
87JtMt74hcBF48SEib4lzTQtOqfs3QF5nnwTcOu+OpuG1Ss7FU6Lanj9OgWSNAAiJ+ChzOlMa/JJ
0/VNAFvTOpXB1TFxCHWJnw3M7Uz7FwhEVQNvyiaoorTC2GKHlQ52tYN082lnJiJETMHnb6qu5asV
LHGNmSbEZiGgS4tyGW6ALgtcS6AP9Kb0nLDA/nIQI5YtHlM1VXlvgYkwglX6kAf7yAfFYVOcS35V
cSDsJ0s3oinBQjVO464O2lMW72js9kLARrkilFYuY4WTGaqxxsstOXSyEm6PkxZTFdSwhOaek3EJ
V7BwY1jcYogprxsR8wv0pba8EvZ45AQctcctny45VHqRHRttaQpoAU1focFNHwoc+tCQQxSMmvwM
ioyMRgG30EJc7RVBj4x0sMU2clpK+bdkW5zPVOdpCSjQ9LRoE1kFuAqfkuho30Cc0R14oH7dK9w+
WyxG8Jvqc/R9qin+9ybQeaZgYWaydIL2o+/DHgY02So5CO53NNszT7OIvVk1qrk64AE1AiEPClsE
bP+Ve3nMBXNswWHnhVb9uqzN8MHBnGpEiNKJreVdAKBGZEpNQ317692zw90GDOlwaFkCOGyF/0qx
5nNBIX+UGqNSz5Bd9aZrS4I4YhcFs8b6P7qofrMx3qfvynAxeU3KIpC5Nejm9uZFASBwPUBRGGiu
0FWPKSH8rbVcoPHLzCsB2N62aY6h1XFRNgZvDVdzWjhNZsLltanIFFGcX89cZLMYwVRXJDVS0v9u
mtbWExfpWdJjDQvWpa/J6P9FceRnC1vyD+tmdW504GkLnR9xRc/ofz6XCracK71tUyNwPXtj4Gh0
JfnZbQsd4UU57WIHGwyoo3w3TKV1P8F7F3yBnc3HNHwblaY4z0eJyA+bBo2OYXhN77VhjdMgv5rQ
OLyxn38MdEganzkFFU4ICccooz2wa5fR2ofh2xEaoZJEHXcYslFCBmJQi4Sa965u2qdfop26t6Ls
6/WjVpM0LDy9qAX/9L8s9t/dkFckC6Q4n9w5BP2yZ3sc5JOZxiq+PdQhYpeS9vRWhUSJF+xEa5Hc
m5sOpBfGlThhq6l3ymdpTAaGa/uNpvtAdw30VdKgFhrho/6XEFedA1yBv7S64VMO7mEMgXzKZMvF
fxcAj6Bpgt96Wxh8BkZQAaxPbJNQSISissJFTPM/u3nZy4kIOca8IOcm+RPuI1h2K5X7H8JjGihK
Mgar+KTGl4CPXOE3gBP2EdNzYe7eHmAYCiBcy4ywZH9f1taoKiiu4EzXiideSPhGDDH+6Fwtv1Az
rGnhcN78iFKPLX6NMMrG+sbsMExRgK7t5YMa+Nk8XdyKZVYPzS6+SxDGxpUeUVsVrl8WWKmB0UU9
ICG/2R+c9TUjcl/FpmQzjXDlB0+8XeLQZWpxpGI7qs/gU4LYSiF7DLFvfL2VfooVs1SEUYHU0Dss
ENyyvB//hfyvv28LpWRtZXZT+QJfefBHm6i/MJlkWB9wj2iOIwHFI28Bh/ZzHe4R7aUCA/VkoBec
jNllsXW4nsgnLeW6Tr+w4zQwtgddtSXqzfJjv+eRViRepDOIC1OVe02daPOSdK4qwhCYEmWh+iFB
XkupSdPjrj5FZqwYsEgapsYKHntMNcw5RSbW8d3uxtsSbs4it/+RpoFBQgep/b/EUYcsu76reh6M
3hR7pC74AmO8XZbDX2Q0aDMjng89lyL5P/0Xi1ST9hXbRxl+oZsT7S3lVMS5WIAw0lnkDeM/q2Q2
6zDl6tMPgdYYx8IkdhrXKzbyHuTUD2hdosdjj4MsAH1MOvAT2bFr4o3cehVrLaGapLyZj4b4BRX8
6OGG74VaM0tIUhYoaQtYIyFBrccOikN+C6s9rfhYXJPX2nKkmULFTbkvQa6+mqdOOsU6vqLXLMMZ
9sIGd8jpl9wljDq5Pj34s2G+pHvlKylH/AHdPMP+anbmJYsWyYUh0D2dOI5jKmupqNsPKBN83anw
p58/4CMMwJ55fjRKNvq/+f2TJ4FA2wLA129tugS8v6fvAp3Wg6j6Aeh3/67fiYHV7wP/LjgnxK73
3scHuIGXtjcFnyiY0m6CPyE3Sbp9xXHjcJUlIJNjEgS/9qbFZRAwDHgaPcN/AEaBQ+9Ef9dXCInw
tmvVP35q38Tjaqy4/hebTI0htmrM9PBiMFJw7OngfvJ0rnMCBtRFjCDwF4YLH0ZuVV+2ThJdR7fR
7zwqIi2gbNc8xK91EgThABwWj+q1vlETvxTIA3yJOQry8duBmObSoeTTSqvwuFfgStDvsau++XNN
TOjVPJ7n9fKLA795Kg9yw0vvocatGeKAxtAjwH4z54CANe918JqreEOK1eoMGkDR3gx23V9a5wtN
lHHB1JS9uSPkMQhBTM1dQ30/feo4yMq4sACseW/XNh7WogrZChYYHipQOzW/PzyZsr+mBofxuaJe
xmE5h94p83ytv4QtlhVj4kukDhmuIqUP3Aqxi6IvFFCZPAZ57EG1PvBf6nXS9m2E1MFKp1+ucw7y
Il6dGiNGoyhD/2e3XuOLnONeEpdzhQ4YJHTOxqZ7KCLe51+ZuT++vu1OgiShT2sMQdDIzYbZsE+S
G4Vp2A9L35PH7FLiSYaGQL2wCxy6iriArhKQ4Kuk65wamWAN7KGJF/f4hn524xMuvdo5sj9HuwRx
ZEDCpxHZOFHphhAlpr9/q0rXb72CzgE9zk1nfKZFkWv02aUEMGCuuG9ysgchykS0VPdaT20WmQdH
pjOGvvj/S7L83qkZJye3kuGChY+O8at3jLIzrCJ5GPuDBFWPkjq2QhCFJbRxt6xeytTEzmUGgnL6
xZPHnTjTXY6C4yiOoiM5ELYfYDGJu7Le+Y41FRWxPkmVKrF9BdqgI4jFf6P/+QHseaH/t6Goi5UR
gYWwfqcRnXSieSJTRlByyTpqalHfynapa4mwHwAnbr+lq09DGC273KdUCG5IXKuRZhHo5l5VvpDK
YE2IwTEXaY/6Tl61pJvRnuZyS0neskdC6SdNcfFywzoqgCRfGk7tvIE1NupTH5ppOy+3gi61WVry
ViKfAhnaPhZQoTT4Fh/pxEi8HvGuaq5b8nUaevBunHSp8EN5AoejK/6liINyD9yK6vHVqrV90V5Z
Yfz/NVrtdjgPv2GdG2mGjLpHKk8XjJWlNlhM5H9uU3YVsjPFBCGaVex/hZpKjNwzUhAM7dad6QLM
lzVJH+lhxsHaO1ynEqsQ/SzmTA5R/9x29Z4kLzsp8G0OUYtri+pk1MtHUdlvPH27BaEQSQHyxf/N
cp40piTNLGDA4yh89Y1a7C0CDT9Q0P8XzhCqcq7LGd2iLQe5+ouYRno8+4mvkMbFzCecoBcwpWRC
l1C+M1i3UZkq+xfQpL770wKWrAs/iOlBG31qIEQnG90VA+tGZjeoWroTGXYPPfZEG5CIqDz2ZRez
jTr4psNrxDXvkkJxFu94w5L62R3CClYe67xzFoyy+Jlzdx9rLep5lFRBFmDNn3u57aiQT6xWBBMs
Bg3aM8aPLWyH/MShTJEzas7YwXgoZPnisowYoS8ounV6Zc1DMBBGYye8Ej3XG/qXvxoJens7hNVn
1rdvfBks0sgrrWC062TmG079fs+cbeKcloiLGPR5hi0IEY0z0K1913QhGK1YxyRgR3fAqWNs1ve1
lt1Vu/jGbKVVxMC+qDaRrYdCIlWFIdI/8LCGm46Or09UwSfskhdd7/ACqKfFHK68ggQWxiIJ5ScA
qkC/BHLZpOVueyLse1lp1kESFuNfbUPnCFw7Qz5Z2toTJohHdquQoM+UF2FiGDaLPUqFM6OXXys6
PPGEfpRB4VGxtYTeFlG1ddY1pG03uxfzK8RTLm5glrHVsL4EWSD1rzskSUSalQJtXOgrVhmxf1M2
oMsNDJGCPsZgJr+wYa6ylHPhlXEjccpRkXmNfTK17MKLlOAsTXXlFfbqfqEyTkBsqpY4BAunNSYC
kTWUvk1IqNQIIuiVvrasuevyizS2+XBJHjLJHgsXeTFB+N+tgPZNlDFbwuZxiUqDSwtm+Irmhqrp
t04034R7avbLfvxaMfDz/2UG23msR8Tr+wqkj8qegC7tfhJ/UIefLAGuJ4zP8DoFY4WFs2kWZ698
SWTp69jeeod91fuVUSukP66akt6vUKqF8jvhYRYM/xuuXowaR/7weCHeHjuV31djjXezKm+6vJ4X
FZb54DMIGRxabdG1FHH4R7C3C+4BUSIJMUCO2jLXKQQwWgjncPTV2WRMZJSazbCKt19KJeRKtdSR
WI/upyOCTFa1EyBiej9Sgk6xBjJvD5wRSdVSzToONGVndY/+lDzkXtnxtJLSbUjQ1bZHFZdre6xu
oh6n5k4xCGqdcG30kLYAmuMDjug++TrlFNNWAN7KN24m8P+Wm9c2VcIVcAC5bj62vsTLjbNGTT8/
BHRWzw384b+vEGbHCftE1/BgAv785c4DmSx3/5BXVWbr8fkp8oHnqMWfQjQ+7r9gSGCbpDmvXIhB
Te89nwOIOfXJ88uVCcA9MNOlptD4ZQ6bz410mdPB0BE2w0BrFne+34iyX5c9BxSsnpdawmBwAWtF
PH7Pbw1ojft6Lz8ijW7fUVY4kBOhjn9wz4EW9EHouq+XE913sU3lx8LIMkPzMSPbseRE005xG/Pp
ccD7EnaMjJ2ZD2T2asI15HThElcnziq0iRHwFv9+SirU/zalkoE9ufEMWDz5RRxQOvxuf2KBooE9
RMIcfEW5+Mm1B7OWo/dhE1K1Y9bfZo8uoh43h9waaLrzGFQ9/+XYmD8lFNL0UnFDCJx3JegmLsT2
EDNqqXqzKZMIfIlk4Nm4AXZi0DTCDF6aUjKUbyAR4GlbgrmLFOhPzwOrXSf+gve4YNXiC2AZ77B2
C5s20FdTGN6NHA/XikthxMPPdM9C23ZtpI7Iv5KrAJdbcCBnkG4zAciAE3xP+LQP9PnkShgN+zEw
TOfkLYmw1xmY675uhGs37hDudH82bDSAnmyKT+NrHDanCrB8l1TKR4qjnc9iDwp2msqqNBJo3HE8
CtrUIhD+7kr7wKXiYhxhANzxm2wh/gle2UnFJaH5GBgh2DNxJF8lble1YWlnT9Q2KppEUYbb5F5H
CROHEKdA25i7x9y+b3aFy9K8UV4EkgUyaXa25rIi++PPOMAoY+wNdVFI06X985KXmNA4hGYR1PLl
AcP38VDGTyCSnH3rokBQpVqMzyrqehtYpTA7KNwLU4eNf9Zr9Z2+xhzmbbR9m+/ItiHx/1F6Qjm5
q+/+lvu3O2cL0BN1JdEWnRE9U8Clbd/CcVpk/5vKkntxMLXJjU2S06RBx5sUQpbpkB5p5IDk5j+n
Okot/xdl6x34VkynLt8JM3bPPCAx4BXVdCgX7gbxMuoJY7yHoe0kF8zt+HYZ/nWlcb3SJLpVl10Z
f6uWDR2rLoTErrMDY2crXaHcU0S8kMXTlnba6LUs6N0Pld+TiZcCemyOJgRUBQMGY4iieDDWz53Y
VULakiuQ4ghGbK5klszg/uB77C5TBc2B4TMPNCjUVeiMEbPZ78NQ+/ASs0Mvd+YFfyFARU3KHY38
Q3kTQ5g3DgVpZwVOIuNrRo/mitVmN//jQl8E3HaX09KtGfdeZ72hOy78OCon7AJIeFK93IfLoPc1
d5zzc/tyQrxfqDCTo37U60ILOERO1bsp7t8QPBktlMbr+e46slN9jDRv9fFgMoBOPLTvRKLmDkXa
4zPw+Jv264DxXOsSxGaDg7DT3S0/D33/upAPog+BqyphZozRkncgqIhC51h4PiSv38nItMYulmuB
P1vj7TLeXQ1jN9yEDA/2vj/hH+NXqt2U88LCErRTZaZold1+Fcb2zKGvV9JQ2cLpctxBlRc/sZ/u
CtY0nwQVbIPVrGQIoktNPI+MpPZ7gaCH/WjJOsN7LEVroWemfs8upEuIfgL5fXGdMemBZXg2uKjA
Hh7tuwMBI2D2YgicmEqDy6oyMBk/sdPSc/MwaNOkU/waCdi3bMlClyzCwTd6q9oeIKfuSnSEKjBO
vK/Mo96vZfcqch2lbgL7saGlDzCX2z4xdmhO4cmE6E3a3vwMgoLUktSnMIWG7sZnm8YyDb/ldAdy
664vzBUivVNtYaXnJEMeXaLVX0dCeGAy9SEfmtd774jdzWWBL/znXljDbfLc3owllXVsr7NnTMc0
YWMF4bhpl6vckvVFV1PSawimIqUVugWuTKIs2MTuiTlebR9M33rmBDZ/8vszMJGcGses6pDziM23
uhqhXPhbfQ3a36E09BH6BZquKDk6MUsfksgv+xHzrvjmvWlX8tj2wcgAzUEryEV98pS5m8seuFTe
wYzbcHWA14kCTpI6MgsN7O2W6fDFkB7onFc4msWX5lNrgN+mlSSa+eJU5qUySDxUv2PjcGQaG46O
+oArrtVzIdPRCkhgsL0mECEEMw2M0ib948o7KJau+uogQAFEsPRmL05zp5ph7K8NIor6S/0jTLXA
ZftSq7tLXlNwuJzNZAnVGI17jBiS5icOZok9uIHrGleyTaC94vGjMLZohYMeH4mHugqfYYrD/XdD
WTE2jWMB7uhOF4ojlAXxNVROxWo/MilBml5JQ7AvoitqGnrad7SCArIIJ8phRrGpORpYeXA8ZUlk
5dxnRzZDjjJSqaBl9i1B7ge/huMHQJSAh1cszAyg8Wb7vy4zvBldCV2IrjwwbbBvRQw/MRVxTxtR
cI5Rw+HWYqSQFuTQLdpe87u0hRic07pPTbCelsINuxh9ZNa2JyIp65OPlYPAku6unDExSL8UFZp4
XiA+WSr3UUlzBzJL2q5VMY4Wps7M5+1v7Frrhr2hDFoW2S0uaIBNBQxhRnoJKL+i/Gh+j/BRxLMR
pWEeBpgLD7TJqLgDRSGWXqsTBbOXUHYugVDZKSwWcgiJLmkfqM2cSWcdMXA55Cj16qmhbQnK8BGL
3yEB6pOu5fIps/IQTQjbtQ4CbqA56csPZ7P+7D4jkwYtUczQ88pay6iiQ7YAlCIA6Po93YdSx/TK
t0M6rcCNCi4QvNFjErq7PXDcjbDqmmfjxtan41iqsokyoQ0vvnF/UKAeh4xOzGxfjeK6V6aYBTb/
Wum02Z0DPyDdELKExB/UzzodjIN4XY9esvHxIRcLCx22LT86u1IZ0rW4D7Wc1xidiI9fJj7kp0Fg
wGf5GwaNmeRzqYQ1ZFxQ+QrfJc+uhZo3dWRGw1lH125eJD59b78D67k7Ek+RgQ64sgLhqwVn1yht
AGndwh2QO2zhxB2cTbAkLqymCzXeyP7oSopBK4/bJ+0o2sndhLqQlAazJftDCRPRsciBccd5cABz
mDom7Asx7e4umWQoAPsC/6F0VT32tR34yVHDM3esquCKWBIgRKghBjag0ItiHPmXyVzcE5QcK578
aqNo+klmK9nkrvrN7a+suGRGzvvLGSrqKk4rZFXMRna65moHPJPFyUdE+iPajnvjHWR8u0uPk1IL
vvGlgFCPLpWtVEzMczhu6gDZ8jNHlCvt7xTmZhfAQRyu48v1oU9fmqi8iwQvKGnwv4In0lVFs8vE
FM2QXzQrk+bEKfmQWVWMwOLo2DAx11x2qJx6HKueD+JTXC9/hfhWhTg5DEZEYiJ4q7uov9uibzm2
twZNnWDHGoC9vpC4Yr1Ur5TST2n+pB5UllJeDLjSCjSOQmTLJ/VHcpJwHvuZSs8WSRRyONW22yIJ
NobD2HPkO16yx9AYUsCr+ZYSYkhZSaSRsCFBIEhHzo58UaddPGxVvd7ORs8+JayCr588HCNXzpnH
j5K5blrHTe+H2ST2E93x/IdusgmJApPWVoZ2OAylmy0SA14B7eSWnLZ59NdM7iTuYmQxw9dO6pcg
Vv1793KbojFXfDSVbfUnSnnqFnFZa9E8vitPkYUwwjlDj0c4qemkFPZiDaiAxRkAu+eZvjJElyhi
veJegEyrtfGmTNakzeXmjfzVhiHNFWa8SsjoB1eDbNCj1Di3P/BIkJpO5f8qtDCnArcp+9/QU31j
V8TMkBj6GnR5cmydvF36W5VEfmo60zhhPIpmMbkZi+mDv+muH1rDd/CvSOOge/qkUweMRxc0B2XX
YL6krGkPd9mCboIPmAcKV0qk+ZPh6TTNGTmSE86UlfVP0KKDd+i1huecef4GGTLBVz4km7EAJVE/
mRvApDTg8nGHZ1Ew3rTeiRWRGRk4tCSwTnJr/oOF3oVhHhoOhkxwPW83cSd74VnzuU9eektYwMct
rY3Ge0HDnjiGLKHfDcyThwQeafBKwU09zOsjpMLceqtVXFU6MSz2P08L5RmttmS6kajEcP0VYR03
I8AShbF2F7i2Yl0ZWTh/1X5B6Y/YHER6F+A4NokrCzxbqRmmoEWKks4b2A3Q9lp5Nxt+6/ozCPfE
S48ZzkaD3lhM0oNS5zOTViWfhp1VALDNzR31Mfn1yHaCoxb8DfcOHRx93w5hGsSiynssblW1dbyQ
7K/uQXAzwkcn7RKTThPLw6MGMK+woDRgOZHKNcFh/Q77X7YEJaRB+G66hvrzk9/FEJi6JbXGpNxP
PN/AFPNnp4OrPOrORKCSoC54hCIMqeRq0LZuRiWd0BNIenvSKStZLgAK+hTZ2YmIqxsBD40mBwxL
oGPtmkf1dPshISYdO6RAk153fmff247jT0lBt+5D0ilZ6STRnNwMdoC851orw+kaXS1kjUQYZxTa
w2Kf4/8ZGLjdEyr1A91WL3T/GDs/sWucVnOi0b6060Ibe7X7vIvqHQrdLTsViHEAXTPSAvwcQSut
MZZdcX24JnBj5egPI6IqumXa7efE8zFeu5zEjq9MLJQ2HZfstyHnwVPTrved8Hw0zGAfbSEGuTxb
wGOhuhhZTBpnbyN1IEGZqThcpizGLa16J9R74kmzDJCKYMCevFo1/lnOmftJui/j/uIhmDdWBiLH
b2JatLT3gpbiVdQGWuV5HWV14dpP+16Cy3yFC00JP5xAsE/1anoMJ9LUq0N3QBcbxWRl8mt9iR8i
rdqDQzQy5tTH+V1JZr62EG8oIydeMmFevcqd/HvzxDk/7xrFk5jofrSPKj+fcZF6rOralKBcYIwf
2rWDV87Wf8l0kpC7i6LnGHpV3UcREYOlnaiI0oGxXBSMHEM7j7kp4LSgGvzOqRVAT4bMpwVxyGs7
P/3GCKzbqYYjtS7MciFLRKz3apXkVzzDaCka/2LeIaAZqyduX47qFAKaeyJ9lA0pNRS+hs5BvyRt
4Zfk9GXaT1I/GDFpVZtEEQWxG51rsZahsGga9+zGuK0a3cHxxPEPpesGSvJTLKsKfj1BwXOotN2u
e5AM9DXwEBV/fsMG7kn43JrpS3s40UK0XlDSFnMGytOviWGgQ7lM89fnAFkBtboaA+UHJVrKyJod
hRM8bEsMuIrfDbeQHZpacTWWRPOcU/9J1e5JWms85cuwQey0F/TumXf3d9xQqZ7jxdMbY4CxLnke
83t1IgbXU2E8cIKoalGhvd7H1H7XTE/LDeuadupC73Q5L3rKWuwgxXwm7u93tufG2TPy0vWzXRWa
zxEeSTi/QNkC0vETZZrL5vix3JGhKsXkQc16maGj8+XBLxWil5mO2a+N4gESo7gQWGCglTlUENKd
uCg1ne3126SCLIawypwFJk/jsp30Zl5LihOp2Io0zCLVkXyNohA2pmsr6sfkN2g5SdPZoUQG9sT+
hVOkS18PMcZZMNiziJ35pBIh/+wTf3vYLsEzu3tOutqBZstIO/C+3pH7gkeDRC4fCXOyVtVqApm6
4e4Jgf4FxlvVQed2Bh6hx5QsTWDw3bIIiI34AMnAZ+6G5bj8SkKhCGTbRCGHhhHOJH10gOyeLXip
3hn2bI/QhpfRQ8iCxfRCQj5bSg2jFXkKrrpp1Xqko/EdAnfthhKljwGqrIxTh0OAn4zBktBMqU11
7rYxyouFW+Q1dIGz3tv6t4RUb02aTQWim9KwFsLpfprhOLEwcjsut/IK5GgxiNgAbTaI8UnmF4If
T4JlSckoPML8IjPxApFUZLTjQat5Qa6Fy7G2A4mmN81/yX5gO92k5FmAJN5/c2mXa+NO027DeK3D
oAX7n+5QwORqCRdmbDc6jf2TD6oKM2KTZPUxQPT8UQoYiABjDRG2iroisOPyyUpEMrxigx44tPcL
OpqgpTRllg6sBDng9c8l+h8w1Hhe6yjMi8cObNTpzK0Op1XMYKwJermMDueO7TC+oMkztnY+Ja//
nllJ3h3bPz4uja4EGNaO6BqNi8jP1B9MYN3KnCQOvHfSg1q+7yhh/Pch9mecvrDHEapg3CYHq6V2
YX0rj9/Gh1k0kR0O7GQeAP5Y1GrmlgYntqRjRY1/idOo7j2LMe3FE2sP1K4uXhzfuv1cHVso1MHC
ctGQNs/Z1N82+Yy5hO+atiWllQwaBd2Na0dKb1h7pHV/Sn6GspPcAMmurYqLWaFschvV/UdpC1ks
1ZQz/hkimotWlrrSzQ6+X3wbZqJd7N5ldyOlOM+9wV99v2SYykX8C+PQAqhSN0PE1+iN9tFPeu9t
zA0jR93kvvxTQuVlf5oMl350aprboX6Ly5H2ZLTRHjl1WY/q5Q7UBpPmE3PDfKfjmLSZj8ktzKgv
ZbPrQnvRBVou2EDcz1OfKFuefwXh1rjq03nya+9s6jhDDQWAI+OezjkZreb3YWA+RFNoS9hV2yQG
4CvDVR+cNYwNCyd8g3B/9MgNz7SXHfu3tlCW65+esDtZy2zVqIcmQpLNkqmYkTOVMYTpA+fR+j5j
k1UbP+WwS4f9nOh9VXBmGjPGCGCXx0CisZ92gxZLqdUafdIpYOumY+XfL1H75TlWNAPnwjMGi5EV
hKuuQxkBDjXtIsgnZ5Su3hFv6hQd0Oxn/6P+gDlr27Nia3509uptdX2n2WP6F5MelJ7FezHpOInX
hjp1ymuL1vKV1Xowm9FN4Yt5v+Jcrf2RyJH8KhpKW/7Rh1Q/nD8S/HBBGGtQ5kILTe50kyKm7oaI
81Wg6PCG7pDeLVyKQPa3yMOrTZ5lbA9D1oa4oWtJ7g+90btqtEM0N5ZLA5e1t6iuB6+ke7Am1yP4
7eAMU2unpVp5Csnue3IJNjm62ylNtelyD0T/hHt6ox3zttUE9lkErXJc5Vj4hHQKXR23KfzL+GCI
0kUJ0+bEQz947t1pmfLKuhiakCgflFcgFKXgGB31u5rghbGWSD/JdOOCmP/ulnFZTeDvp2LKTAR3
oost56aSKx7Zcs9bO7qGHAjUUQl1C9jiHo2cWHSmkmKkfowzZ+eCK6MszjBfX1MSPCaCoUhZMjHM
tpCOPE2LN3PFV2Yrr2X0GpHzIXbsuX8p733scXo3J0LBAmLRnVaQZld3sL8wdzyTmNdKBqbmsDDb
hp6OQxlyQC4XJscIUoWlM4/109JjHIudMY36Jd71exDeYzXjnLEUu4B7xggpnL5A5wV0t+EIDX88
N4CJYXl3OYxkKBfnFC37xUOEr+l9DU0KnTh06vBG6YreVpC+XQ5qDQhK40HmgEkkgQV9MBySxIxh
XOG9mOrTY5UA5QyLsX3wj8A5FsV+Dm20/zx03+AeFUrrxpR5oPfk4wvtvmMdt6WLiNj9ZnFpFv9+
3W33fUyx8p6z4BTwHifFzOCHrHkAuWbYGFw+u5C3v0O97rdQtjlpoeTskRGM72myc6dowhT9/wBr
m5mRTxlRDHPx4UuZHb30HcTJqWfOHa5/lMm3wACQztjmAS3nbTcloZF0uIKUNs62NsFefBwdgVaR
m1J3ehPYF1W3vGceX7ReQb1jj69+nt1drft06wSd2HBIw0ELF1xFPLrLRYNHa8Y2LNjti7/e2J4+
jSMvfjY6648oQPlaZJc+zL9HWJIyWFQyL3/70UVXJ1Lckg1CTgno1bN4ZaTy2EWeJvWUhHAe6+s/
j67wBCVYAqhe1ErhTK73JCoqs+ItRfTHMHIiYPNSKUMSoTSbLoP8DnLICcVbEf9cytWKWFukY7Jw
RiBA2vp1usoEdW5jGPgDEwXGL00ibeqRL4FO3Doj6uqhPdozXHLhzcJboTIZYXwKmeYVJahrtfGT
DO/3n3E0Ej/iIwvOjHCQ0FpqGUlgoBBm0ijaHmKuYgaj0cRtgMJ3z2k3L5l96y6XqUS9g3qYF4c5
U7xCF2YuHa1DbEDejWWhYdiJno36AzPbundmHFqnh33xYgVkiThkH2C479SQFrXIPkZGp9S9LXbz
kOX7vOfC+8N9zKAO6C3TwV4G6CuKrTCDnfBzayGv/QCCvmuRT86J1F4nl/Phzof5E/ofRtb3pa/7
02BfKD7SsZFVO/H5UDuVnq5k3QEeQbiavywct9/FWp/eV4XBsOqpcbturNgxqvrrIO+Hl/xSnwh+
E1C9H7hGnYbTC8/AqcS06X6tm3fdPL85wSmCBOirVOG/ByLSYekwmfSUHZRq+fwFCBYhOULFtX4j
mTGaN41QAu0bt9r7o2bAVW+eJKQpR+c2LpTKdD9AgTWEV40P3aWLYLh9AYbBMr9wPhRxLoL9FTXy
lLrJTQ3PJmlUSrQmqFVFLVpwbKjrnkuLymSn98/NDglTAIRT15n4E22osAF1QGg1kr45LqLyH3/t
dpSIl1BoJY5asILYHHi1uqiNE0OH2UnrHimd5BLfUAHW00vbszkTxY0+aM1Ul2iHCeld5bzWl/Dx
EH+1nGYp4S0vSF4p61iWWIXOY2IpoDMYlXS17cHm/2nErUEAK10tZrUUYNc7k1orDCzqdaVK+R8P
9jkzNjgHXoTQWUr3PsksAbkUgRD6pEVzdLurMi8N28uoAmnJqa9vKIMSoWfzRa6cTEk0dhmKb0wr
7eRW3aglp1rpiAeBiFXdeHO4Fy3JJAl9NYMVj+YzLx0Qqz0HtU1+ZdQ+fUac3l4ZTGDuAHIc0Fzo
J1uhZ3CQSgTnAfxdW+Quea6upUBRC65qfbOghYejblNtbKmJO9TW9Rt8S+GRaPStwv3Dnrc6Gl1z
HhYNXSEJnP5ejYv9Tf55MXE4HT6eh632V+k5Ms1LIm91ELtjHgSg0TwaOMympVcvpqzzIfQP+1cJ
7Q720+2YOW0eLaDCyAR3e6iZ3gG/+z3riSMrGF4l3kktpSa9g0Drqa8oMbwijqWXWF6hk5n/rhAQ
qHaxfQp8bCsDxWZ0ruZq3VFF1YIZiIzZVXS/3d1n0BzrxIe27I/l4RqHfzrjbmVVDzjIi8Vsq68I
KqGaQwl66bwujefqXh/hxlV90LAu9QSp1EDFJstc+9KeP9Sennb+mwKevhrYiFD31Qzu/cLr+0Ei
P12tEgOb3yeNt/rFgw0BsdK+WncpMsNd/bs4VZKN6hwKtm1vPo8FvjlquerLxJkxPih4UcJug8AU
zx9H24VTdXMT6vHC1imbaOrxC3p+KbNTt8BBL2lKpjXviym6Q5r5wyRWrvKLHioO5WVztyWDUIYi
76RRxk9/qKZfYeVnPKHdJiCF4UKEp//4O3UAavNaeec+qgpuvxYRnVMdc9C8okE1oJrH7va2IkCd
ARFMnbZh6Gw6Ag6tn5V59N7j8qi4pNKNhl1TxSqYitdv5hz97BZSdUJa70TgQsJiE736BIBCN6S9
5Fr54Dy4R9ugLE7gp4M3V7ysI4pQDpVDWXjhULkgImpV4CPXVtl32+eXUGOBRa67KHlLd2e+NIgJ
L8YPCE4SDnKaEpgVs6Vz7KdnqirNyYBBVqzV5RhUnsAcs8SR5qaLOZ3NIDsS6LkbxXtHxjPE2oDL
XhdExB59rTRQk6CtV/ophxH12UJ55v2bWgNzC1FJBOVOyb9Q/GecP7GLURnM4Dtx2pAbq+UEXnCy
xbODrxcUC09MYt989VwaxNyXlxN2YCv/ogr16ISs7/qowQKVwVpkBIgTkCC98Mv9dmSEQM0LxxsX
KO65lr1Zoux/TPiX1HbkS/RCoOB9sd5Wg85eajpcSCmoPtnvpm3FMdD3cqgfRAedSXAjIQ8UMe1p
/b7gM589YtmcWdAr3GpuLST/lPT15zkFZMovLYw9hs81hz/C3JiMZqk53zlW2kjUuFo4mU7w2J1h
zHBpXvuHypd5YvE/defAa8R3hGMPqjLLSbNwPetnxlOgeXw/FvLhARMflsI3g/0vchOGgm9+r1jo
TTEiQf2h40ilt4Ol4oyGDmerFJKD87+WQhvYsFyye9EnZaD05qcd5lZMwlh5uI0QsTrtUNYklvhr
+G7sD8clKofpNr4YCmeS2NjJQ9HXJzBBWfJ2KA3oD09CEplgx+b4Fi9LYdamyHaHg1Yq4GWbx8ac
M1PffibTxdHfbTjh82DS44GbkUh1vSZZuzpH9WEQGhgIF3+zNtlEOsYf6cOrSR7IyNJ9CUqDWooK
rH7yj8OPOxG0Cco5YwAnxTRy/XvJ9c7vYTjLMyp1istEGCa+R9HL6duNBCH9To8SWGFdTywew/Kc
qwi7e53glEys4p9tAxW8WG6ky5jGpLnXSF8C6/bd269eQiVtfh33pkqgzel0lAkPsn0U8pczgwyi
WT3ta0Gscvpy3dOupv43o78sq+KQmE1VCRJ+0vLMIrKbnWBnyIMtlzqZ40fPLMEtjYmhEZd04Y8+
tgu23OjhUNM/aAOtGcAPohult8vVj0qsS30NGrAjidSwITJXSN8XWro5KOAr36tsHdxSPbSgPhVf
QssL0RY6dr/eJo1ae18fpo4lS3otFaHBcsizUhbJkrQ8VrZzXgIrOR7ZNBcWQxtEQCB+1N7jfx8u
HkwkzDYZgoC0qADRDzA/bNl1vjfEh4q/QHZmNYVzIIYXiwhYfBXQBGyM2MiITEyjB8V4TeUw/ctk
F93UhSw+RA9b/svJ16xhqCG9yWCDzUP1gl7Z9oqGLp9ewvmlvA4dLuD2EyF/2q0el6BbFa14IHxW
+fh5L6rl+M8YCbmWIib4ZgDzWHyr5HWZLl1eYynL/Zq6t6jY13gJzdA2CiVd7XtXc6lAlN/3jpOW
hVfyxbo+Hbv4E3UvZRy5W+ejBKHmJ2fJl1Ze68GnTGoSpHbfuLjp6iKLeZq1xFa0bRIKYzS9iqWB
s06T9AdtdasxeAbE8MGMN3jg367yBYh1VXxmWHUc0tCnRl7jB+vHGFKISeq815gh4uY6hO7GH9Cn
2GZoki7x9k2+WniBXAWscb5qq3ZbcgQ35UN9sfjcsA6SweTDZsmgWIBqvG95tOaGaYtwbQOa/Hjb
kYMiMwPEvfL7+7xPUvN5NCbPn2cYzCRjW7kNknuMIlz+P0mo9OM79f90sFFowWQWt75DpHyJp15o
lzLfdDlzzGzqJWOQL0JxnKycQL/FGUar6YBFLEKCTLlPEYFRWx2cmYdzyCmJ2OB/UJ/hPuEFA77i
JUHnjnpayvM/et60AN4RW4h4I4Jfa1pX1CZ1WQ1eyAAhvwOe/mIJOBewuM/a+0R1ZlABC45+vOjV
R9F5LLSsL+i8LEcqNlrtgk+HmpdzjDDElPwmPjxqJd5p5HkyoEoEZ+WJFUT33xfSYJjGZGOjaEPx
7NzPt6Lmp2S8w8duysbdXF7QYJG0H5cRrYdLBaIFaA28C2KDNI6L2glzTuSBxCgBsLaIQlGoXb9+
XdK7ueKUS41UseRz9RNF4YMmN0i3qbsA1OjxI6QjX2awd9x7PFIUL80XRR0TVYb4lWXjs0WHOCiu
4zeeVPqa1TFyAEnyvw8igWH2rnXHGJwL4kWkMUCb+49aVTY9WKvGtW80dkVTKLdOd5hvJ2jydiim
mwu18dZXdPzYylwsrdmV3dJRXVl+p+WEzlrHWKd/9qDZDldo/IDUJzldKtmEyhD9iSl4+F/MvhlG
5L7oJ5YVtH0Fzp2J9jCSaE7w4oOjyjZOQKkeJ/G/kcG7sztwmMR552/2JkOgwhVB5mWyGoXyUPvm
FafN3MrQGS01yq167MEZJAoAUqneeep2ahgc9s2VN+9d9BGNeK4afHDu7UBkt3T3ar0M89DKZ9J7
zyTA/VD3I01xOT6tOAVCrz3+YtOTAl+gCe09MeWjCIvAU90AqqEId8H6M9O5xaVgVuEyih1C2dwO
ZuakSdcCD0qjEhKv/R+NRGreqj38UCW3UHUYJ3XuFDnnPt0MjshQZvre2pdi6BaJB2BK+Eys3uIQ
A3k8AJ54bTtX+OOvU2dqEg2/eohBlxSt3L1telyrKo6JRdm0hST0VyvyQn1+tEXPhTKiZtag6iPN
taN6v829VjTQJaQtqfyxfI05tL3g/a/7vSm2gskpqKldp0QxBfsvKmYpPZZYzECXOEg3E+5RnO2W
IcyiWqHx2DWj4n/ZYVoMylr/4ERfOqDWxYGs/dfx3sorc/+qrJjlEXOL3oRdWSaG9OohdcvxJlMc
qbTyG0RLT3c+VZUWZTsUUD4l1RKvtyQsSac7rKUgQ7MjIAF+RIXmnqMrlM+OdPXgvLJs6HdAhyv/
rhZtLyz/03StQeO07G7u8xa5J7S7ixlQbxHPD1WWWn6aci1p9+lxsUNUUZY+aWqz/QAjIQ6+/V3+
0n3ZTXBb49VA+dLFCltkBnMRdJqhKuwDufMBAxJoiHNyWdjkgyFE6iLaDxfDXa0zgkzqVmcC8bTg
f9PWtfjBx2ejGZz9Y2ciTL4unYaJV8zY/5JCpwNXAoQ4q3gy0xYJxW4jgID1PaWz1kAuNKrP6NPP
Q76N6gqWfwcSpmdJ20gm9eZBoWp4DIGZCCShBdv+YVkqzvQOasikTW9X/0tC8yNckaHnXhLLBKL8
0O0Ejq2+tWd+eJGh7BWqEpHF3+fPiSyqs+/jOLl/rj6TO/jyI7cSczdx7VyvgGolYHdfLcjF0y/r
4tBMw5IfRMtkI8AW5JIkDaL1GiR+zpy8+q80OIFHi6kL1QGy3QveuQAzDvxBmxVbcBl7WFuQ7eCM
XWM/B1By2n8fLr4cESQhsJ04vYwbxTbHsadr8LcWmegtsvsfHVXvtZupO7buxZ1R2OZb+Vfwv2Fm
sPbkavGZwxn9Xk3golc2zZW0dAhj08OAQXsColNX5eyxET4NRT+4p++/a2pESE9EDzz+p2ETodWa
IFBf8fh+xHsd7Slm0mP/1LCXjml54AueiV4lesHGckJsCgN5hJMffrWshIlMaJUU1hUzU4sLxU9Y
jIKZ9ooRHuLyBoxets4X11sLR+gNUd4i4nZlDw/D4sMvAdx8g/Rr331Kr2wRo4uQ16dUPk1CiTsG
rpRrUbNBf8LkKE2KS8WNrfkXEFLX8KjZ2UH1x8t+9n2us+Gz/3xx3Sw+qVvdkuLz5biPALrWyjfT
YcUi7Ff13xSn/sJqpepyj2XFd7AK31FNskaNjouFxu7yROHzRbXTsY949SUuuROaNS4UpsL0n9qW
L6ggSB1UrIqGECWEtPSjwx3yDlXJA44Q+L+WpWoTiuKVlElh4dNp1XQJUlOJzK/Tnnje6ISSOCOD
og1PBtRnsXwRtd//DkmvOhhj3Flui15I50F48fF5S8EV2hd4V0P9lUoR79UCJ0ksc3x+gei4dmJd
SKiTos0DGoN2h9WWSwRpB2vKkd0MLN5QIbJ5bb7rySnZXxCG0WjoBI70rTR5RZwxsU33dEqQB0Cw
3985NWZDHX7MrlV0DmsfKFXBURm4Ue6esLIbWilK6ZpVBlAnXyOSB349cDRTN2CZWKWTgg0RqL7m
YabGgylxLsvBShsd+Y4GtWgRXeJ0ADRQ764OfDQO8mPu97zEw13grVQaAOQBcINrLtw2AsJLCg0a
/Tpf0/XhgisTyzWrwLBuXIspFNUay4nFspulsAApuKxReE8lE4X9jTUtlQiUzDMS7A5fuyI0tFVx
XGv2eHAsPkdbLRZ2aTJp6dPX6uUY7OVftK6YGIVafLIjS95klSplWrVqbGtYbyJvH2fJgYtWvwQ/
Mbg4kOZe1g2D4SZc1a91yzc+UjGczGYdCWgnQI//3JrZyUROnmW2f+yW1sxyXh9n/xhEG8bNHsSY
67h5xzJmTfO0m2LhzBcB86LDelOekIbWCfkPRrZct1Kz/qUJ95BJ+Onc5FycHLd49U25wQ079jNy
DNQQkwTK05oLnZNDZIg7yIR0Z8rakOvDkfADgbq5u2zpXVxMuEbENtHDaf5M9LLsN1o/gmDHP6Uu
6dqwu4tueqlWlI0fqoId8kmSBA1vqLRsaeZKYWnSsmiAjC4NKHw4jRsGq1qm6uA1ry9Nz9iGvgec
9V9LO8RGexw1yDQFe3x/Ux/tCyU89nFOj6VkGt7CVBivg2YrNK+irFTPlydEvEQH0jmi/Xd7Tsfk
Zqk+Qo9euxrUB2qnAPTsjxlJn4huf28G/GENRMhRCZaSfAXzW7c2h9N3nFu3Pwas/iWEgqB7d584
1vq2XKD20ooMiXvqhJORMxGhBGPRfTqTkZ991Ebz2pb1ZQUNStmk7CuWacvxftdd1L456G+erTvD
KSwJax9D+6RIU8AZ4NTRUyp3EO3rnNz7n5ehac6EueICooLFwVlFLatOVwO61GG/4qbGgiSNtaUS
8JFK+65Z8pqDZanyUkpj7ilRU3AUW4VNgvwRP9hUo4VZq7d6he5fn/Y3iKbN2PF4kXrZ1fA83Rwo
tn0Wzm8BNY3ZQlCFJCZdyML7sRNIh5Y7venwDJMDrHQX7pzMO3E9XiW2RIb92udKm7PA9qseP+en
3//oNbPRVcGv/0HWPeFNxDpfsRrj2Wmj9d5gDRWdWbUlvJqZpmBFqUtSNh0NfnIheoVC1LM2HbWb
v43h5Rfkg19ue/ztdxYOt7NL9MABLW73UVUX7RVXHWOlmgvW1KuiyhvZl4hvlDNX2XnJmxgvCmM8
/rzat/UUWEHeKxKim/gRS6Q71P8+xZzO/Ke6UU7F9gHdaId/kBiWM7SqwqRRZR4ioBS2raVpUKv0
AZPsESLiEh+vxrzl7Y9npvQbfS7vYDAiZycP2/M2oP0GYvCBg8I4jJlxRZvWKwEEXCPsrV98RbHi
fPQSDwxmlStE2TRp7Idi9BdbYlRpxlii1AstIPpJJgOHYR7nhOALVre6U5STro88iYsZ9H1u4zVD
ccMztJg3sFWg0Jvrcdu458VAAJEYjG495fYME0TH6riGZ9VuqUksaKfv0CIwor+6AjS8R1uvK+y6
hlP47KHOJU457r1vsm1BQpoHcinIM1LNCIWgbGs7T4cJfmLfg78oJbXYZJedxMh3+4GclGGr/mX1
W7XR+Tme4YDnx3xe5hQhYXSdGMG4krL9rdnslgw6eyJkc7uoEnwoMaNTnbZJ375Za/4+XnL2hHLK
ec2qiSXadsefovmKHtSxtFk7VbH1gQaZKFZ1ZXk23dsnpnFI1NqtIyLHpMu+SN4Dtse3c3EmgwDn
RxCswVlYqynqwi/GfMEQptw7OrJH1of6ysrhqIko2W36Ht6yjzhbYO2qGk2jRX9cSBTCTSDQm/IG
R5WvfPuc7gm3aSOGswxRxUzmd8a8S8IFvCLa4Q4A8TSv+jm1hwwU+u+lzVrJoRYIRwJLsY0Jla5I
oMM7gkXRxxdLlUN1xN4caN7e8Bc9veb14VPe1ViMGlO0pbU9jdM2oWWxvS4dYqn7mzXmUCB3J4hm
NEaxf7IAOS9VCsEoXXRCDlugfh0vQfYpStk0XkEqXlLH7iuWyyGcGIE3kOxphBsKkzqUIKvpHG34
REn5FhdKIhdFnq5qRumFL9gDsAgXpDTJSLSICOXtjO/M2WQaU8oACSF2M1AFaShTp4SFou8M0X6E
p0mZRD9te91bkS0Tl+BxpsgGK+8qYX65OJHO3rOHO0fGuiru/gt3emwTkUCndEf/V+KcxT7jh6Ii
HLXR6vKqsZLXC0WQ+3NJp/aqzsOoyeR6u3rWn8M4ntOyntz1cX8keB6a/fVQ1qp9QB7VjcI6Kiur
I5/P+EoTg8T6IjsKJrnd3ttalJfvqvzJ/tKoDfH3o407jzAtLsT/oZcywUAOMoZCzPOXEzw81qAV
Kt37oAPoRKg7JqF5qDJsSOSDLb3oE8SqDKjfbKatILXFuYhNLT7A9MiHpyGTZdiH65+PYT7WeuQl
lzu5pWHGoVtqHiHwU15C3E1+dOATBGbjOHIA0u+2Pr7ZbLo6H32izepIqnAAQwz4MOQuLpISobpP
bqS7T4PNHCCRF5d8ObsfXIBtiYYwnJq2lAPRlYBf/3erCSRgb9+0g4IgHQDZRfNGHlajbELDiKet
htm9dy2pVR9UlVAeEWDZfaapqy8jTN5x6KyjPfjmYUD3Qe39Z3kpCeufbwHP99799B7JkTGEDo3T
8D1y4QluzJt2PttTOwXQ8BzQr9cuz9PcIHWlU+Mda/biRoTn3PCYWIYboedADI4VM1ywUeeUB7bu
tRRn50hF3FJQ5GYZFk8il7Nz7+mOrIKNhnRNoldE2CuU/0aF5C3TTNgaojjvOFBkYSaJkp6u+vEE
ezlxcF/xIJ1CLIcX1bpT0aPyyCOD7/MfBfSKYQZ8WrliqAWmAwVsRBo9AewjAqum1t1Tl6BKqWfR
lolNSMNqm0sFjWulKkh91FIC5QMWQ0GMl9xiB4bmk6CZsRm5WRUntQzbx0VbsjcB+YJop+sYi5lT
kfN4mBpUE+pfLxr5TPozn6tsq/yFQXPqLZl5lYrH8EFypMOnqWN8/j3fCy+RatnI9Co22XiGbFCZ
f53c7NBWzLDZuZOOtLt8h/L5UH5/Y7TTYPGxKRyWPxxjpimjGSfwVYIRSswQRsTOLF9jv7vhU+sE
VQaN0x+GPwmB4N1iVINt5beCLz9ZPrKjYLz9L/J3rDR4o6YebDemQwbwyXngbjOObLmQFZDR74uL
KOBRGouH6McRdd6hZ2lezMQSNRWGpugxOWYidXQa59DTeOPa+69Nmu9fShdNBycrtUw5U59G5bhZ
YBI/otpEE8YyLKfFtXd5Vv/E1IFXlVt2HNqYtyGA2Jx/PSolfPzzA8+N5aUmIhVDiuSldGCVCDGP
crdhgXS2SKmJV3KiB3JAum5Jvj0cbkqi8WjzCu4w6DLhArooB2dmoJwAa1MRe6foxdjYs8tWlk4E
L45XzLzEBHw1909VF2YqzWOPPLtMn9/pxkikrA/AuspL/ldGuS/gE8tjl2GQ8kguAQG8N1stHKzt
Pi6bkBoHUmjnzBUpJDmhDv+BKLPh6h2N7174Ax0l0aZfD+ZNRBt9gXoODlQ5Z0PYKD2o18lxCzCX
TvANJNx1RshauLa9xCnCIxVdeqfZB0vMU3VDs34Q1NUTi+cJfqCwzy4DpG/eXmEuLgXQ+JhpQDXP
XoWczLlzenMPiCJdH/2A900OO/7uKhIcdxuNNQM5Yiy6hGuv8Uq4fYdDMJ2wfDXedTNQ0pIQMpsz
opdqK5I3mukE8IP5kod4/ejoRIa1iCOwvp21jDMiT576HPSLNidtjENc/pRdDxbhWmqp7T93nx4d
brxVKI1Zsl9Oxn6ZH1htsfszglC1Qh8OO3brft+4pZDvvcrH/PupF61gTaMibFllCZZ/L6CM/faj
zlqQekkx5B/jvUReY/pa0YF5Of4LrCFROfwBQuro2lflJz+Ph+eink6dud62TKlW9G6YWsdCoeww
Zr2B5unLd3cU2ddN2ho8C9gDmbcuprUPRV2hGyHqpS7fpXybyGLZjGVEFuFw0AV3F1OXeGBko7x3
wNny3aQfN4u9vH+s2P65av31i+aeZVSIzkgaqflXlVOwz1l2jlE7xYtao2LkrM7UNlE0XB4gDV2n
Q8f3cFraJrwXD1eFo4hSmPwxAwAgVJX6B0qJSAC0KNdvlBtHYC+YhlVDorrRfs9SoCNQueuLEiEF
zHqdiKL8Lel6qcnNEftHEpNu7SgpNhOsiLPT/33Ol9s2rOI0eDoSnmU4Z5MUhIUlDOnoQ6ZEyo/o
deAwLv8dA4YAp/LYXJ9ZwrgPQnDr1W9BepY9N5IfZZq1rlOxyPU13fMKXFm/IJLhLm6hRJGCDH88
dzMDh656vQJDMeYcjnEvi+vsVUNc7iYkLz7evOD1d3t28L3GPN7kefzQuEFhAtKZvSNPJZJjG79M
PypdNCF7zHSBs1hMP6OxfMftZM/1/ByWHZ47Zr7pINOhWB9YZ2c7wjeGpaBokQ2sPwcd/LM8pEWx
zGu8DDQ5yqqKshvoJgHWmwdgyjvnMyPgt/MFllF6JPWtsw+gJ+DIGk+i9TCMtov+3NV40E/TkcLI
LR04ekIiqziRJDXsCaC7ljm2qLbBr0WS6HBGw2Pm9NxDLThun/Kb4q5uKJLcbqqIf2yblxfPBlRJ
I2zoY8lvqdAKKOol3ZAjlOnVVLB3JzI7HRNZuxn1T+U2LRd9d1Zgm/lqtzxWCuAcdX3bL/sdoBvQ
6G1ogJeSVMMcxgFdsAWuTIWBSytgoUiTSFxkCU8nE0l3XH6azQj9N2YExsTUZOZCMkrPJpaFwxOe
hgg83tseGaIjprujO+MIW6vyin5ESrfV3ta+dn0RA+/wrZPrxFRX6NZvpjoMGjx2Dhy+dyJPcgIs
BDRPEX88syB2POstNqUTfjZAcO7nsIZVf5GIiWy+hx7nPyj6Nsi+rQxpvT0v8wlFBlBwifRfx9lx
mauUFObW9B4RPZ2LnMwLPuSZNUlzvuEsqHcXRCCasgRVqvy7GbPgk9m5gduA7czayc04MYiV0iMn
YvgOPM07FaBZbEyfiFJqVXBhSj4nGRFvMwMGTkTDZsaGhSyRGjiyLGidfSrHzI1ek/W9tCXn32C2
FqTsqN4TTxCbWcODd+SdWMpY2gGw2+8ueYj2baHazJzgd5alhYuYoXUHiLMjL4McyPBShDaTPjBR
LJMYvg2M3g+qT0/5TtAV7/6r/Yw0RdiuWz2sEneP9hkENlZnZvvmgiZIZdCgG8ZO0G2+FsY0JPnP
2lyypjkbNQli/jpGwvv3Ycmm9KjGmqDnXhMiRWpeceO4Rovdntv/VGToGGD5SI66EyrVo0dSdrrB
q497L1wn5Qa8SBUHvlKg0CNM+I/IJEeWcypKR+MGErKmaDDvgp9aA15PrBUis0FcyoSoVGdmvq4N
3a86MgrDQBqOO1wNMEMqp+2Fo6Bvj15+AiBV71cs5/NQ421IVmKatik76NRnuSsb2u2d1A1tMfrL
a1uWg59oQS9NOKGf65qLIQbvhv7HVUKu/S8UkcIIi/Z3qmAo9zihdJneHBj/wtja2IvU43wKRgze
jNlBqha/hq+KUmKvRuMjQF8qXfKqz5HbWzy3xz4RTYl5B5uOcXBwtHOcGVlGTox0jsQfL6W3Qk30
rV/U5OVL1Lqbcvlm5XuXQQiT5WMoeYhJ/gdE/dadZAv0ksNSTqKmj95nnYqvq0zZQLTuJP2ri2s/
GYpZ4fBqwB+ySZm43Bdpng/Q/m/bxV5ZZOlEMRH1Vmg1nMcSPYAzLqpRK/l3Ch5XO8RjMyU/INrB
rjrC+7Oh7JrQ/IRt9dt9mdHoOVn9Ks6ZNdMaedbHugLafCkzq1trXNzHzK4MhWKQyCOxFFrZR+bf
cm9I/bZFf3J9hi0qDUXx6jvES1kfxyvGZY/5Q3Eqvro3ECPvE64Ak4nwM/9dha/ICp77q/FOO0H/
npdg9OiMMiQ7TZVy9gX26A4va0tFFelwe6RAHHTRFku1ShjQ8+hj8y03Jgo5E0SuwqPryXz643tL
3R79CPJ9cRvdR9dNA5lmsk2A03I86bbnSxBgy1cgWnriBnVK5NPf70hiFtrjPaU26xoR14/3r5pe
9sX0ZlMuhzSzL13HHNNkpdYTV0Bu7YZlsdysXE+z2XklkuxGg9QuMEjSkCLHr9lhWzSQuqw9s9zC
Ix12q8uWrXKBFswD45OwJSI3bNQJBBfEcuyQJymmJ03DIshT9BmnuMnWl/OAheAqihhIcwxADojA
v0P+ZbOv99pZ33A/Y3+bAzsUmJtUbfwwjkCmVbkTNqfPPwnKa89v6PSq7pxorWGSEulYYX1oP6K7
WRylGJ9cWu5cRN7CI5jG51TRSHb56m6fgCbUBYVopG8NQW9pncNcxs3LnXC5IYphAAcc1kaSF3AA
LoXkGmIla1vSFjaOVmn8t7NdupB84zsYEvE4gWgeouVLPJcx4jIgCXmIu4Do+CXHHFEwyGAi2Ite
Bna54cw2dSpZmeLCGypluV9cr3i5sgo7tTPXRVIMQ87pJXobzjRH7QZtHME76QxfBAHPyI35fdW3
LRwLgcroojbbaybw5jHuPU5Rwjzf4+G+ofLgFyxhQUzcwh5G2BAqkMHbH8lH7oyBzT25W67qFwMp
/8q7blKCUr+PqFJDdE3JOf1EtTEZj0jlkznLM733FLwYXYOYKaQ3EvzJ23edaxAzLIGaZGmOWbH+
Q4hMOGHMK2qkCkys4pohjC7xfUGpRIh2zxZkThyq+wDPYdGpq4uQ7cOvb5ARYMg+2xUpjOOq/r14
HAj0ujAcz9GBFqt4xsw724coj5dejgWjhlLaU5hP2/HsSc807YBy4zanlPLxrMn5Lv8GYtQFwHyA
4ek8l6hNU442Wusw74anNt/rXEZfQmHzYIBPec/EApV5M3USAqWlZraY/UupLl3Q44oE9EbCdXTN
930bgV+wOLAOle1JnCAqgTi0VcMRp8ME0KKiL9a3kcTVyYBjWTQNGhHa/HqRb+kV7buz+zwVGccM
ccEbS49e1KNsfPENekZN6KH+gqVoxw5kmKUpE3z+OTYyL9lzMVNvpNcTn3KSFdpTW46Yu1pnHH9i
CQTUS7183MlWj1Nz4N5RynjrUJzfkG7P7yf4IFupHfMJYvDX5Qk1GMdKm8pjGifkzhBrIzcPg90A
//6SBy7JfvGQG4NZV1VDDrNkod8aK64u4PVo9evqQzrgxcdL6SyE7IHfKpEo7VnvqHWj2OZj8ojJ
1QN7Jgp1VILE2GFKLN4fFQNhTjHnzNMZTSuDMzw+iHOvkjTcudmbWT7THhT63okHN4+jMgIFz+Qq
7kmomIHhXeApwE6OaJ5vgucv5mV0H42LfetfoWokwJBiZR+ltTWlgclcvMa0isTXx0iQOfm40oXQ
3UecXZrfW+tU5hXQ7V4X/DF9sY+JuOjXBir9cg0Njl5zN0qVooKCjosoqEIRdnNIuu77OxeZpuYF
2k+TDVdoAU/CpjjdkcPG60eOFbQWQQab/6RSJWH1ivuh45IJrhrbRcpmMRXCoxM/NERX2f1GVIwE
M6BIaNFW24Emf4yAPynbbRwQu+zsTaZWOxH+HJWeZLoJZDJpOc+FKjoM8FxdHxxJVMzMIWnK2IRT
RMoEnUgDYU52pHA6caTdfKne4Qrtw2KLH+H3iMfwbP+2XKqfXTP9hxcnqz6UzcYtG7BO3ALNGdhZ
UbrzIZuwCJxZ8lDoio/XM1W55IouLAyhfrfp6R9Ot2CfVh2TuvMav+UjAxq3wzCq95npxUadqG5z
UWkmdAZjAa85sc+QcKwcEv+GF05aU3dZoBXli8Y7qG2rpu2XiFssEqtCrMlOMAxSxVs3TCbrwhqD
IQ+sIs+zsAjnG+CKOcyDqeqWdhnsAsIYfv+26S2X8klv8xE1rPNm6jFNYJjqVBUz1ELUwGt2ChC7
x7LRX8V9cH+AmewR+pqkdpolgMzJdTcU7HPaJd9DMWP/+8x8EVbUI6nYPE6UfIWxvMf2gERmWfOU
CZQluRX1a/iVh7SyXuj0THRNZpCVV5BhNLWJRFSUvYz611JsZDeiKTVL4Plqx9EpmT4adL/k/Aoz
bLPyZJqaHl29Dg4h12jMZKKblwlIAr7JCXeyPpX5tPUEb/yhIlDc6ta3EHuz0qecbuAbXwb/LsUG
5olyuLoRtph3LJD0qSXLDe/96sZMERG+T60nlbE2m9ZP+/SPqcTkm9t43LP3dbPsV1bp537EC4n6
OmH47MnpmoH4hYQuoHo4cKePioNrVu6L80WNkNG4cPXDzLHojNdwcH6YktbPRp0eRLqHu5WWWrNQ
BRvQytaXNDGpNoBB+tW68yFT/BfCVeyD8C9TBnuHNaPZl+mUiJGXZzAwafIz2kVoQAeQPAl6GMo/
SXEYvsvYaBnVP51hVo8b8H4J4Wstl+S4h9w4Z80P0QBGTMhUsZPprSpH5rrvtJCQMNkWIX7aYoE7
ZrAyLqs2QWr6pOLlUPj0yEFEteb5P8qtChBHuBIHCFikCi6b8TrBg67qFgxtm5gDskPuM/jsZl4Q
iw0uEpVGNrtDN6DUOXhWxewJb0M3uU/ZwYz5RFBCy+pSyoqW82/GtakI0HPkg7FH83wWYbgeLvd9
Gxc7Upvn6kMgWgnhAgdpi8mX96gukjK23N9GTeozuyvR4pBpbqvLfDV4acmkUXtbXKzlTMvKusnp
cTxOhhMnyhIGEuhKN7lL/RVEz76E98MpaypJijnUturSPNmyDIFyZqtAqj9Uu7j+0Ant3IiRYnkj
8OZnzIMx1IXj9YeEGmKkLHCktTpNJoDAT2SKc9KUgYOsiygoWC1jVj0GQ1gHUASHVs9O3m6Y2upY
FmAZp+tjeVyZtcWh8ozv/8cRv8DtBsarxKv+FZVjnOxwkQpkbZcmPz5NlO3/uatXc2coDv6nnj+C
k3yDScU7hKOTsTD546kJdFcHhnrElzhlxPlAve3560+RAV5cysitdNpkJrnHtOoSDBgK42ErZDSF
3sGJZWb35HsyCLa7VBB7vZ+A429Lo1PkeMI8GVXxhP70welk6AcvuQ2p4WckfbzJYcLLakgPxoVz
oOID9bHCrq0zA9CFcxFEm7Vn139cLwYD+ljcbhvjbxogzKwbtI8KW6wHkfjSq4Vgx8lg5iZD8Rxq
5vEZ6mgwGMwQWj0RYpEHyTSzQJLWr7fk1XCnQ1qiKpIuwVJwjUPOOI2GNDJPOYltW5LTTXIuTgPG
l+PF7DkvMB4XlVWPNEYvk8HEeX46ohNZOVF8DffCBNYGlh1XlzPJ/9qX8OaGhTHAtLszbu11HeVM
CNhZ3eG8LqXfSPLYiBaMQAGhsiSHfEl3k879cccMJHHOW9vrEvyiC/r19Sx8CPSrJz7AwAqFyuEV
wSXTmvmSu/ztnW07g70BS2QAlyCzAcQeVqVV5sIDDlRMzQ8sDiWMHnY6w2QlDB1EBTRoXzRi1Wm+
8rTzc7BZuv+F8IIcKOq85lGrJYKWItnRcDQnfYXPNpGhXEAZimz0l8a3Z1VwORwPEanelspXYk0G
DhmuXI7V8hVwq9i+0mNAgzVDDIHhxj7YeLMSfodDpwRva2H7AJ4mWq8XWhPmqwidbk27ZvNA7+fS
EbtlqD5PW/xjr8nIPfjD26j+kZwqttMcwV408BYC0w+76b3wgpkWFygHF+Bidxjgr9H0oOlVOA2A
fUCYAHprvlxwhJzWHiMThDU/w4r2TSY43JR8q/5XT6qMrG7hyIQcgsmlmekCJXrZqSFiAv2aXRCx
jzTMW7ZxNyuODVfNdr3WATtxtIbcHWi4pipQ2lwubOAOytDt2jXk9VrSx4fQAbNzke/cQbQ1vIRL
4bwER1cYRa6eSkan0TTOy8b91TQfAs4OzUQKLOnbgsvnxENwjviLmAkTPEYwwKkh5J+e74soX1xr
AAj7bEqiThX/PNQBMLpWR++vUk6DgSdhCZ6cW960MZ5l/SZhm+idM1lT2C5H88BlOdDpNAkCJj9t
4oxVJ4Fabc/LPVstISYgHM9AkuFmR9HdAfxF5par14pfkwuoE1AM3KRhai/RxtO5fY8uh1lBQfHV
kJgHoWbD6i6NA0tYRk2LAy8KBPEXaRWQDON92SHKWh8jmpjea0hvbbE8tDF3VqS0kp93M5/Hh71R
7j7mbwvojnWSL2EkwEKJSqGfNMxLj7SiKWGNghEyB5Wcv+RqAbSZ245GcxDLCSW8tXAjnGFPWJyv
nYh5C97NRZmUpM/v5LZW7/TTUt68WuzqVqFt+wCbDNn4sD1wJQ2ZdIUh92T667MOxPmIcGT5tPg6
NDnmqifWbv+dPvpw2Eu7rYitpoMHZ9P6bl2GJiLZzSaETgDy/nURlIwBwWkiDzRKOFqzWr1q225V
I/5vhuzQq1qhT0fw2+PXa2F2g4/jgvlch7drKXKEI/xmh9tyPoJfQAt7xKH8sEefh5woEauzlQC9
IoGroHgmQNBqdcz8xTg3vjZkqCs7joRZHXuALufjAhhaegQEi0RcvbuW2c7dnZyiJe0LLSOwboEE
kn91mpI2o6++YXFkBlx7HcYjh+asgOrD8PFsMXFos5RNUeBCaihvtobINwfoApYUpi9BHLHs5XtC
CYcjNbde/CmyIq2BI+8/vZi0v6RUzJ2f0qEUtuNEefNNnqQPWh799ftFDWYgo8lE74ggqNLiXsfj
74kg5kaZZG7+Yxd6x/1RIuXuO5lvHGpbTWLHoQu7UgNBdwM8Sz3x7vGeitXwyQptbx82ZmSkOcQa
tuBRa8Q/3dqCHua3M8O8juLOX0x4qEi2Us1pBE6c+kmZ+lBl8gVGx90wbTg6RGWS4xLzpwQQnhOt
jBfw5O6/iMlIVd07I2/egNesCu6NIgPiU/IKS4cc1ahMwja0/QEv1yJrPDnKu5sxUFgnvVbO+WrC
xAyvEGMlzgi59E9asZod1F5gqQ7qZ+++ZDXtgw/++KYzurPQx8CsymIgVyS3BEs2AXE2xZbH0wjy
1bGK4kS108SZdoNeY40eYpxZEa3g5LR1gkgbZuvoHn8jrk2mjKfKWyfy3RP0nlk2+l7WDoIBupk/
8mi0e6pbsNZFIHUBizzyVOaEZaGzcwKVFTyTNcy6crcGXgPuj2XnkSUWTmLJxkX56sj+5sPOWhhE
PkX8xH5Z6z+PCaNr5gDDfaEUOJSQlyKVX76Vf29HNBZxFZjhiw/+RmIZxLceF+L5NXHTUlQ/AG6A
KznxpUkwbosA/XeUzSAhXVBlzndRrLjT42XLZFOXXaXoh7943MtMEbcOaPu7bohAQLfSLdfs29es
Ggngxs6pMBjtqU8QZ4AO474eB0swzpsV+ITXJxyzHhiE71gefNWtK9VAv0yRoZ8ih2EyGSB3081G
mZTijjXSftfp7Mw0Omom/VVvBb00J/InV1t+PgU1LtgG52FAnZZXHAAwAtYtbiToAr52tEbhfAzH
sIDVEJe7Y4Lt/nnflR+PAu8MRamejZjBSmK2Q7V1UeFN6Fse2VFyJIap5baljZgJFkIckCJ0B+Jb
TYgnlK5pQZg8N8NgJcySA5e2c5tEhQJ5JRjlA+q1Ttv70YT3VIqVX3MntddLAGZo6QfQ0JA1KnJk
yS643kvCnfvtg8c1ufBASX5nLu5YENYJUeGY0tKsVDjIx4be9JSxf7tAiE3l5bES+/TmsG7TILw/
PjU1VfItVrPO193qv/OU+q01WS4up+f3/YuvG2wx06joBApgKleVg6ItsBe4J5rH0eYNSROmmSVu
Xl5EBzfaq9W6xvnxzPcc+NKJEqd9eK7cD6dVRucyApgeJXRSogaJExgGLMXQuxf3ITv5z0TRg8Oo
QVTG4I1ukqpS0aqiq8D79dazvAdTou2vnq3FLRM5rFEU7BOYGizgMpig0ZA91b7ge06EnDIdGEkR
lih05pOErjCyEaxRIxNaOjHQWrZDPazTBFOZmWcuXQSEynP4+5IaCadFAD7Q5vY0G2mo1m7DDFj9
kYBGb3pYBP+qLWXAY6lySG33SrN/YPesrSl/ubZ3TVCwhkoRMr85gP+e+yNpTbagXB4bp1NKdEEr
T1IanHVwRiTsTkSv7Te1imsg/KTYi1zOGpQZRpn89qjgAB9mDBTwJaBNiSfL0zzu2CLn7sE4gR6R
v251SxYgAFSLHBzkUG05aKovVXEb6rW5NzXyRs9qQm0fDkmAFpPCldPr0g4KngZ60ia+1ewD+a5j
yCAvMaGlqA93einh5zJPiaJ3F8d+U67W5bhgiGj8+Qg2pD9DhmMgm5RTepaJNy0XuuSnWPuNP2oJ
eakyPf20fRzVfh65/PHVBw/1zLimizPdcqmihuKrUoj0kIGGMdVq4DYoh6rWfIyjXMH0VmK5sotS
Uc5yvy/sN45XRWk2oLjYruxqWopK9AQkrYvVgYsR16wCMJAKXLi6VCvPc4jKWEp/5bX1Sl0T+Uw7
AnWqaCz9tJiE1986J85h39ZCgpQUKPA0WpF24f7P2Nmop7E1CCeJaQSDWXfenFybTi8d62J8MxRs
mq9qWhzuHHk9PPKttO91JkWqbGSnizFj7cIsQKqmobMoG6yDB6ulzJm37LFiKbJJ72CPAEHOdi4G
Sw/r8CeWlUhOZ9D0XN4+LUSAU6y4zgKFmvfBIozVL07Ax9DmFgELujN5Lo9PxSuzK0WDDYfVSJgj
1CbAH70MAwbPvVvWiS4UB9cVivXqUOs1UGDTe4Y6O0HqU9wIgXBQqYDuWtNC8/StikbqytQFKvBc
u2nbNwbFCpsKHR2wA8wDz2pHljEkGfIlWzpIy88AhTRHMDG9xF8pxY9C4N6QudU7UCKZ8tkZg95q
0+8HWImkhBxBohKV2n3PElms/6u9A2jqoBUJhi6u9ocDCcdbDE4h/1ITKY2o7U729QjYReStFQML
W6WSdgapz0UzkvmK2rpBe58vpxs0D//WZpjfTVwjV2/qCxbTWlt6Z47+b+yv4j8/55IddomkQfs1
Pkulphb706veHhC43gIuvetBN2YLEv60m5lz6DCSPhlWNDtMkvMNwF/pSb6C7R3J57cCZDr3RibK
ngA8dsIensFg1KU6e3Is/a16Sa1AvbZp+maTCgneQUi6x81i9qoAGyfYLKOfdKTyig3Lp2TzxP3w
9Gu+GqQuEVK1Ojxl2PsTMkPtOfvtxQ75nYsRjbGaYJQFZ5FcKu2M5+fJ6JSSO5b3RplCOY4TOddY
pbHLrqtVOltgHqH9lTdsdT4J/TXPNpnSkD6A3brC5vBocvFEcvmDsVOvTNPXDXYzLk9bZC4cRelh
u1g02noa1ywms1HOXlZZlYTyJ5Q0d+iybPhaZH3iOqNAhg6wLFhxu+avj33YeF1fWva9ewBMmc3Y
YJnkf6n6Qa8GWDiGW/W5fXnHldGBuYTa4ueDl+4auE1z62YuJ0xT484GNorcKE8u05rQNZFsgtos
pxO8bUsqOl9MQiEIalId+ZhgiyWlAKHIioOHVsRrxKqndEIihyGnO+Ks+T9cyN5LimeG6/yaOYy6
huODUAQ4FpMDxgjoUtauTMuDdz3iYhWIhYNzdPDd0Koqi1mxlzrxIBNK+Y/qtZs1mnVIwyMx3ttj
cfeMo65lWQvQSPJB6NprzwnIOrbu2Jy+aDoViRSQKBOm9+Kzw17Qm0T4gktmkB9jhQU/NUQPpw/s
SOgI7gYlGS+5eTikEFvrszL4YTzBw6I9g8YfUgZgTUcUHEXbqBTUr9SYIE491bz9oIfUlwhHy3oU
fc30ZN8G58njfVGvC01XMBBbId7GgGVcsVFINAEajtZH1DeEZ24xr64FcgVyR3b+/Qb79Cl4Hg3d
4zUDh9TX254bRIWTiFkfIVKGx1WjOf4mE9jJ+OMHzxzB5p2P1QOBknmQ8wNeSyNnSrR3wrvv6vcK
S5yyUkWmo4XV5UG3PYZsG23USqX0KlZhikWZ6Wcz64pNMUD5qFgU+05VHLyxCaM5S4L/A/Jgl5KH
nj9GNWUzuAptO/dTnAu86Mep6WfAjdpGVjOfbP3783lyduke7uddLldAs1BYWXXxd6Gq3S40iulA
nIKt24C9PKxZHtyxV+3dXGe3mWvDvd2vWPNL8Di91glaEz+eH+7nvrnwhASXzhP6pdWSx5pgf99+
CqN2jskCIsCkwqtd5fTUCZTXDZEaA1spvPHTPxnQ8o6ZA8Wx0ncSXPOw9Lm6fRO61q4B6v3qxugG
kTelXTOvD3fdQpZuNOFHTmDw6eFJqTbRtLRaMuFNYMCanL7szc7nsnVqR70yBgpAtdPJvhEake/4
JHOxLy+g/dj4uUdPyjctuo8Jzwl2uKpfryzW9L8w1Q1mP6iZoPzOlDH/4AFmHJF2IzjXexagvRkp
p0HeokiK+Z/vtN8qdox5AnuPNLWgu1BtZM1BkNdsmMO51qifJ6PMNMZYKo1F66FqBlx3cgNvR8SM
TIrF7rYrlFrsgIfl9XKYrBcq7/tHk1YlMiXG9BEcHVWYGOWyoINgfh+nVV2YWDpmYB3LdHbVO5Im
rotI8GPt3epprj8y0m87RmTJK+lk/QWHn+Yohh503DSF+pN0SZo3lKL8mbzsRKB3mv06ceDQEcl8
S2TlYW+ai4OqugdEuDbLXkJLHOTne46WsJaF0b66aWZ7+FXPzVzaNULe+S7aahhzpVSqTWqIl0OX
Xwug7yVl9x1OOrY4ehGH7BtxGlt85XbHvp67S4++bxnAfwnhBP3Aw09kyUvTryYh1ob2IOlfjpN8
y7t1xEXIAwiHLQmz1WqAkXHG5cK/YoaX+83R9/YvzRpnODY4IpP030s6K/Usmz3u+bkThAjMfhbQ
nXNlsno6bGyD4uVosPBzIpMWmNcq7x33jRE7c+Sq0L91u7sNc8xyphmSKIwtOZ5lLx/YC8gGuWft
twx09K5p2zyWnnhC6CGrDRE9cpeQ/XhHRa1b2uo4MrKqoMMZDyzSXrZkwOiqzjdba+ZkvSAwe2kU
rwXmmJ10QFCzq0x1OVHTFBqAfnQ5ssBz3H5aMPXn+TOA3f3/sEt88NZyPmTbBEVs1OmFkF/GAtC9
DCPiCPP4i8h9lQeDssB23e9/n9nfKNE9x1h2Uxznh0nAPCpOeMJsf3fOkaU6R+o5x3Z5ElQiuHXq
7XRGqxtwrxHuVGR6FKBESEJ/qKAlxAPGsGWmY6tLccvC+6CsFVtj3hciVCcY6WLQ42Bb5ZqWOGuT
CcDUtZdzyRqsqlWwq8o96AWrUkqWwVr6bGGIAr7d/ZvNdpQcb6+/tTJqm848tAZ9AmjYRZff2bQf
bPya39s+NCVOyzoc/5KTHmgSm6OeIpGRVYrjs3GK4anHgtteO83qD5Hhklda2tTqygezbZ5MoJOz
2fyPpFT6/mQ3Dpf7E8KsaHeJLjpPINaDQC8xd1FxaiAXhvSezcNgEVxUolWBHtlmviKxIO64exr8
fZtowxOHTlmYlyGAV4ObgsFRf5eZ9QD+zTxvE4A8u6uVCbSKpUiuUVm/9FlsHBfmNFEYUqvHRAAT
N5te0zh9dRfw6R1Y3+ibzkEYX7+Ybtg0Bjik6zc1yA56bkXoVKK2bToSLok5RrwiX/57A+/Le2K2
TMkPM43749NnpfP1JxRAITQhon1g0g0XNsCCW09tXuhYIJRx13FnolneY1sPcE+yzY3jMg8A/3su
WAt/aqYWCKekICMhX8e3eSjrM8xB2o5HjL9MvOmMxeqGqvaW7gV/IinHgin7p7OlN97GYHzgjUvV
y8gsRqaD8oSc7cyAEB8arGdNQLvTvzrJ5x4YX9dTf/8VjTWhwNc+aqMc5oi+Xi7eA0jZNtLQjKP1
Wrjs52VKgkQqgVgmOtnNlOS1nImlrpcfPapEw855fbdPfH+CexHMz/IBeJMQtlzo2PJahX4vO2dK
dz8lfbEyohL+5Jq6K3nXpZwQclJt3nPMjHHMAeVdzztve7VLayztRLygP0fIHRex5lfxSD5ZlOPr
bI9afl+PrgigM4mEnhl46ooxUclS5fI2Z6eK5+41enkXjHbvDh6/orfsm3bbhfadKcoJAshZktWK
dy5ck5KCcMVS+qH+JqXTMNIeqbHcyGsEfJrnD33hIY4QjrBB9Cow1O8GiNRswr0pu6l1kRIUeTgK
Vk6lpnAhjsLEeUuLmJU/55Vat6KZJwXcajpemXMokx9jWwy117695ZFpVfmSMV7hi9m+80SDxMxn
kavJ/a4tLrQYvZycC9qV49WJIg+aUSuSLmFLZPQbcINdasgfWCDSEKF25ebsMCudhHbAV40doaDA
JSzZRvvZcjfB0e2IF19vTVeJI7SBjtHTx2zSNyDdmMBFI+lkN5Wx4c3ZqOumJ6FEkve0GrpsMrq7
Yupue8FXYt9HDGhbkXXgcA/H2XkJ8UnvZZc/8clzq3PHW99emOoeN1cJiIeQJw5K1NFvSo8CyMpJ
N9LuGppfIhCDtHp3LVFnEDljatYgTfoyiuE8VrYpk8VJKQDq8YSJSdW3N3U2bH7Q38vpl2tue8J6
r1k1dtXsDJ6oSCl8guDsWEoydbh3TJZ7mFtEvTG15m/wpMgcL2IwK9JTB7WX/uJ8TbQ91pa5SehF
vlsYqJrSa8Wx5t6qBEqcayQn97h2euwfRdbsNyr3IVinrErX+qGXMgswmF7nFf8Kz6vtleYd84Z/
6m49sGnU1X4eF/tS7TUW8naTgWbVr835AB7lFw8IwLvUGKyjO/lSkWM7yLzGfzR0EjKwvQST8Y1W
taI4eJs+NWgmug3IcRLqJ5OfnkQF710xDR+2z5yCXxqzEARiOsk61n3hwhJ5h8xBqMijRyZ8DiDr
Qji/0+FeUybnodQGx41fEe2/EiNg9dIlnokF/ldgg25fEvyE94tjeOKGURe4wptnHMVEII8/Ekd6
6Y4r+VLfg1BhVo/8EtpdrBFQqU6hFDRxksVl8RMkxV/XQEUZiOof55YhuOPSlQMX7iGq8LXSLy94
H+8zq18QcTXhrSFyJhsPfvsvBpR6J5EOPMnBLiuHLA+FRPCmMms0Y/3PCYyCOsepgF5RsOTfxmGD
F3mQo2f0bJHxYDqaITNZByKpfktbtr4uSEUeFeiAvf+DmybCAO/pS+sdUOrs2ZbnmMSUGgFY6ZOK
Xs8Bgzif276a7406msRcnr6OEOKMDLlUEEYUWi4zheUJ5dBNX2XncND83cRWrrJ7gutcmr3YEFS5
QEe15tdZEWWFd7srjrjmILLwactOBsKmD5yQKFO1ddLZSJJ1v7BA2lRGGkvAYwxmwU0SHtWiIO5C
+jf/fQuIE1n2znIUNqoLWq5iDAypwP7Z09592H8Wiutuoikc/imuMYdW9f6heFt8UExMGEis3Bm+
x5omO30Mx3SY+ASfkjaVwr0Y72mREujR/A6QUnYNndY9oYE5q8eVbvKg5124O32NGn4d64KGeEDG
qYNrFkD+tAu/8H61QSIs8oficmNIIW57tkx6Pp2mxFR+mm5nqS7+9TpEa84p6c/1m+Irhbufxt8y
awrXViVkRiN4Jx7pQv7KeN8B6GEfEexXr2EondmSu9Ewf+uX2IMaOe+JUmbJN1/Tk6Rs3UAztpjr
Du/cUjwZWTViYNXWQePNfgU9yxax1hsD8n4IEwxu0epScSk1H+Zole8WtJdLA6NRGEtdsqffhpIy
BtMSdXLKwvwf+c9AEiTAxpth/2YGn2V0PSbSqqegwXV6IfGJANeA8AnTP1vVSdTBW+YHSO8aP5ct
tDSXixNc2D7RRY3GLiZyQtKrZcGXIMK0/5Cpqu9mumcGWmfGgJZ907/OQuxj5iQj1trIzRGCfvgO
S2/re/m8xibgBoI0/P2l8CIE7DOr0BzxokfS4bT7scWvQFVdQP/k3GRief3vVQWXKrgIvtOjwTXM
HdB9Gy3af3UVEqdVoQyARPcwQ42qI6KSKhuutyAfh4B6kHM7u1ZD6TL7irooEOcHrKAmYDY+rPVj
GHqe9AuE9ZHCpl6XE66aP6+d64BKIduObHy1EriXpKoU7UiiSUds3XioZyng2fVOatWC/4WDXAXl
jCvM14+PyKQZ5y+2NiICHnQsOEaX5GzMMkY56ioSKwsz4eK+RgLamMCfsIpF7zTPclSBEFZ0DJfr
Dh3Z1ZBzmIeVHafuXPh6o9Vvg+0MMgO5bQ31kWTmKbX8lu8Gu+yUPPVabuUlXt+Xl+VWfiaw2i2v
xi/h30iuihCiwsfSzBDrlBh9TrvdYcKS1EIw5EYD5XkpTz4Digl+0I4zXhnUoNpEYZkldcBelhhf
UdQrb7QZuPLKIlQX0tenWCeOZjxtoGdztkgauulx2TLTrgS+KYwz08+2+fj5sIgi9UIfVzLzat7i
3+8qbtmMUbZpI69ZIzhXUP2VvPEbdgos96D0ejdG/Qmd8tUhMb24sRC+ODpgGtLKdctRp59r1yRE
2Ca796peIQBW6zjzQYvTpbts9rNF8FLBuBwYMyOAqUjUmXDM6RLvPo22+Xg9XOb6BOpvwe0SsZiP
sJUcf4Ux+3iSqe5mg34Msa4/lSLvv4MfokqDv0XgYcRtKXCRyKMuMHoykaAeySGJel568d6yy/+r
TAWQHAB0r/8Gmb3dqT4kCPUfwFU0EFUx1UhK5ha6QOHxhCe2lya6oOD4j7P1hpF+nfpHhivByGID
LzB/iHQ/pETovToWAYkpbm6dCW2AIKSLqaB5x0wmpWsuj65oWqI+RMkC2Z5WXXs2ex0WmOFlDEas
mA87IyWmf+wmcJAE6yYbD+0eUIP8hN+aZOOWZ7YqnlgRYkTyL5g2v3UyKwGJQZAlz9nLjdCDMcVs
LxdnuiR5FRbfX2D5gNiSspiJg7/LH2bvR/NGwXcWpV6yXR9LWN4PV8QcARlUJJpfNMX7iu3TnV2L
8kWH36f2iLODaz2tTa5WTt8AtNwd+h/7LgEPJfCwO8/MAPQbWzIDhgL2YMMljOE4EtEGAOgRJ019
fkoekoLF/++Sa/gmYic89YFpDKrBHSruyzUDGVPhYdsyE8VhyRu2k7iafwf0uzIStldNYrNEk5BV
vpOrvG5bz5MA3L3c7iqwdMpWVBOYRCYXDaDVhcFALwYMySI2X6W1uOXb0Rud8V5qnzzuj2HFXcTC
hnY75Fx4dA/LTiXjxl5EwxbyfCAzNeeU4Wxd/+PuJkECYu0iFQfrtVooOaBGKXaSRHVPIv7gwb8u
3GxA7gHASl8UNd6rLCfffBSV7dPAb8uaHjIduFQgj9kpps8uO5GQusf7Q0xAMvRs4XlrD8pdvh+C
OHukQ1hh242Yv/sSRngkov0qKN7tpyEze03eYZ3O2/MLW/YuBlNbakNRvnEBIlz5SaUFZV0iE6nW
Al3isPe6M3XC29Ir2wi54iWmN0eohf3sev2E2jLDclwg2cdqiQ0ChTeLzFj2g7TV3cBCgsPsDVdp
b4oLOcHlwJD0e8cMABT5nJTarjLrf5UcZwkyhk84I1iA1KvU3qtEir8U8DqM2lcpI7bKtqlbPcCg
6R2tV5rGLk825dBp/wd26lICmylQtqk8npd+bNtp/PA0vKuxNrsefQ7by+yvfk++1UTLxyYng9Zu
PxWBJkzwzPBk5xl+kr2ayzpNrAw6WY01JtQt+2SaDf8BNZcjrfCw7x43PXoruXzDuu/tuvYnxgYm
66RhFo8B8aKOjXjBHK0Gy4nSJS3n4xPsLOATDdQNuhBuCeB5jpcyMVvyRbXRf0CvSs+gPVTHDLhb
6pxisMS3tLC4emhwFbEkdWGegfUgni98cm2Oe1Gc6KodEuGzA+h9d4F1D1KpT8weyLkoxs0oTujD
IUm03rGXatl9LUL4ByYNhrBjjjPvNMUQBS9NsEEC4ypCyDLsX7/yteUfMHjP+ZW4wJU6X+hrkGDK
+1lrRJui0uLYPP2Gw++IeInwzocafYmqKyHcS3n1UO60mc6T20n2CfUbBciTTRb/x2VMzdYWcslz
cbyVIV+laf9Mo486YpJHm+oz3C2EAydfshNIIcMGyjNeaTKkSjop0CZWzzDSp3ScZLZ/UZxaW0UN
97PCgLpKETE+pvz2ZKRgUUH/YFqwu3pSlHllY7DgDUOVu7vAVh8NpnxC7xEXcDWgdeCb8SIxjImF
g23vPgS5EdIJXGqkVyTMy4ABU/6LRnbHGmqkLtFvlpYaTtcp97K0YkHUPucV0BwQvpdH3SygaoEq
R71KdQ9xOpaF3IWuqoivfr+8ON+M7dHuzwG1XoPS8xMak9IsSjdbngciv1NYRuVMjtIUEpN7zGk+
EHNAxswoNhFfgbcXxCHG4i+6pJW52X6eoehB+klZ7qIpxE9QAYTYya3JuGJ0zosoOH/LQKovO65Z
iTgQV0oE2VG89F4nf1V5eMqe+DN32l9ojjCpWSD+ceLnyENVeTpTuDKGyrgFpTZu7KYSy6/mqbOe
RcoaBL9p7zTrTEYyzfECHXoAV1W2YCtC8l1VST8S2LjgfwpdvTs1VjdLRlKYyJwCqj3C3nPb5kEd
5cB6jnSW+V8AjVOkRFwgBYetWLJke34ZXqiSq2xaCmhUuHsiYgyqmQZsyUGXFCmyKDIqOdxmu4Ic
0TI+PCOLzRfw0bLErHOU+Xf7BnM+T1dppXwNNwBRX5qInWQ5Go7xauSjmoDWknk69iOuQHIVgJPw
ZXrSMglMWRuW5oxM1Wd0F2xrJVkAXySV8w8eQe2ooEPOhsNrc07NV7gvxK2gi0EeMpf9utDbdunR
cNA0/AslfX91bitmidEmWskb/qHIP75wDfFUldZJg88vivKDBWTYdMFcUCYYnpE6UlabqLeAHe8Q
P0CgLY+cEe4yq0u74jBfp6eBTA6EQrbr3saP9YvG/JSUkPLH/si/rFKmwgaF8tIT9trjkEb/IxNX
SpnHw+F9scJp6NMjtcvYY/U/mbn8LGL/tsgySn2UtePQXcJxtGl8Itjzvr8fheUrU+MF5CkmonW9
BF2do8zwo79DhlMbMxLgTR4DRMUiJzsekFDNPgeXPryqXcWhDA4HguUIjYVx6481A4IfrSUj6P72
qOOVbqC6LgYqc38mVfZyJMgYzs9USH8sldcLRVQB5aIuEsRqUawOQu0CoT+q7BwKl8ZMiI9UgpID
000ZEsqkpkbQrqbRBrVtkqwnn91We12S9tBAQpC7bazVan+XGiwmdarmrgH6WjYAHeodadWzxJpZ
DorUBSXrBMXXUnlt4gGm2QvRsdiRrkKzLP8jEoivwu0rq1Nio6YwTa02Q533kvWrwrknsNewahGW
BJRxwElbq5+BPcR0CyMThT2Js3ZjbIK7Kgyr3F+rSLV32t3IIIT+04qf4rUZexmm7+GMnL275iYD
Qgfgg9aV+H3uP9MbJSweSxw1Kr+RTucYDbiBedSRNzdr+Z2g88GDOZtDUmbd46y7Iw8+DMSI5Rj1
/yYRWlxCM3IIo12s5eCDTdbVPHMwKIHDgewLupkK3GMnJ2GOyZJpy6km8iGSprGUdVsxkVfcUwvR
gluY5AaOJLIVoLvPbvIA8LvaPulrbtQZlvYDquocdGc+lTeIgjFjxYjHYK5EKRyUvYWERUm+uKnD
IMDt8tCYc9kPX8yHIPaoqUK0t42QBuESz3VSFAwxJN4GOay5shcL5HunI0tjWpu+0WaVmv870J5A
QdAfAG4F6F1RKqzlyWVGSRXZbc571VEQ6TpAm3+k0uoiwiY+MbtA73MPnnOgQXERNZqXJxJzmzlG
JSlUqKpcvntvPdt8qOPpUT9ug6zcbk3ynoXhyMtOOjHDcuvbci1lZt+Nr9hXkcoOUNeWUNq9XPyP
vrDelKD2wYoe30bNm1Gkmb59Nsfd9abs8FISZmzx1mqNElWwfYavJxO1dOUmrQsPf5DD5uShREz/
i7WKFTq3y/4rjl7UlK6UkYkiOCglUYhiz3Jae4yF1TsP++dJPQr6oXbQvRKE2svrGfTRr5juMrGn
M3i2JSz8zS9wy7AZiN2Ul8B5DnT1M8ADm64FjnCnUjqxLgfcI1kzhUwRhOU2UMWTW4TL/HQZSj+h
mXfUIGHYtsp0NApwMfLkoQfJohP6He+z82nh4JuibUr+c58J+q6IrZZG3F6gVKzoTB3vrxpcMA9Z
8816bdGXQ1MLvyQ1n9Z3JTQCoE2F014eyskVTWmA6pLqJJYMJvr2m5cc4Li5tiwsyeVTwV7JXMIv
JAAcKl0TlH1V8wdWsrKklsSqG4wtljcH70cy/MjexI0iDfjJmlCaPgVzOYAt64KIiwbEkrTMnP9N
bSXJo/EJqC/kUMgcIosdCPSzGbVRLQn/QQUBTdM+qGW3kQuiaOQfaZXsoHFqsgW5QvWHT//34r+b
yBiEp6b892x7W7yauoc/dk+pDAEVKH8eK++6PWEgl4SQByH+q3EiPH/1iCHIU1dNWkyWMO2xGQY1
P3vBv6KUAtcQNAUUKZ58pA7qJu1oCEaqzeKuMiPuiRPt9tT0qmrnUEyqyG3qvksj7tgyV6xPXIs9
QsvPDT1HTIxaLa5k9S9MkhyOnU8M0G+9nu+oPpWqs+9Cc1494GiB+FAmp61ghpTPzQVB0PoHjnzb
Otfryx5Kkyjtm1YxIXaod8fGsvQcoCAGqKLfCwS4GVOWdyNjyKYpBKvcFMaahgsYP2ilbvOrcZwg
Qqf0GvXZbkcWC4fv3AkmCbkwBqbo0HLI/9M0YJZ+p2uHQL9vuVAvL0Fu3Qkcj0S7o/XHqqLaSiIZ
viyiydBnWcU1eDCiL6it1+6QAkQQJBtOt8+HJRvGJvB4XNFCCUwZC51gryySyD4vB5L0xnsyv7Pm
mqHDjLX48btS5sXW4o3m+449wN2uyKrDJ1oWyuAo7yPCIKmuAKlVrC2JGG9yXVAghF9UzfY7gw6p
A3hmg5SAl5r8TFcIR3BpVPMHKYW9ZM1hyp3EnqkY6IQo/9O0wwzS8eaMSntyTRgpXuceQ461XZsx
/jBdrySlPUTbjU8wwFMMMt3sIfkrfQANCSEQiU2KknE738b30U8ZgIsntuRwXrLN/TG8YPyLxcPl
B0Hq22kQb7WdjmHHcHivfiGQdfEanKp0R0UlTPDSk97DXEvzlpUKI2diMCUnbk0y1fECeg1wTNsr
Gp0JQ/XbWrNTfVjebED+eE43Wp9Pz5F8TGmlrbCBE/CS2LSjvKehQ1Lx0etgLGnm9P2V5XExlX8x
V34axpUQLE0JjSXDFtI81lJP5CcOdqiv5TzdqIvjccWNwwhSP2XgAqhnlBdAPLXnV6a6c8FYI/gC
4oPvQ55vx1ogIYgZB2wifAyOcEo80+xXpz64pPAFFwswgMoWIyByd42GFc65KwA7reDmV3sLA9Qa
dl2OHwUVhT8be/sHZ+ibbE1aQe6V4OGxovgP1uLTz5UbBnxgk/o/69RKSRlB6abTAX69n0SxTjxT
e8IvrmK8Zb9Py6O4jXd8/4qAdctUbXlzoQeeYKTlgqa/JCWl3q1jsOVs8Sglah+BUjOqb83r7T8j
1f2fHQYbllseavIHXijjI0dZc/2A0/mOPpZzPrBqRYqoanugv5jecAC2JTGFGZ//z6RAfs0NiBGB
FMclq5hNYhF0FnvytMFipUOwM0ZUiymvzTWSsu5IxJeiQccWDPffSuOC/8O8+s1yc7mb4lejOjyc
CSZROLbUV0oE8doErbEq0OO3LuAPCEHWuVpwASCEmrZMIGfDOVFGEEMotLZQ4lfAhXiUkm6DkOMf
nSSAJbQ1H1rFVNz47kUrHmP5ucGUUt8F8WJCx7+HsIzt7p+ESu+UsKNMnbMqxt/sIzL1pU89GRuX
z14oqEfE7ykmJ76GMWPFVPtBbrKvf1OXTdlTru+3rUpyADcizp5RCcKyq1ewm7I99t1FXJojKIdy
NGpo7SF0cnGQ21snOVZIpcKPD6aJBSdfwgs+apUwKGCeR65/SCV/CCC28HTgFZgQw0S5GF+TV47N
eAuUyM6Lle+Px3vPhScFynZ61zHsnopWPcdtyyKg0vbshChe+ZbLsK1WCHDylMhmG+qM+Smp4wtu
VUEW/e+Alfla9l3b1Gc3FnqisvF9JEfLr7OmVZUCAd/msc/ZmgbcOTit/g/fxsecnQ4vLEyBwSwx
npTFNfoCfHwqdDse9qFWVYWSkt6BqVVBHuLCg1ClWsW7+SuIAZt/kkMW9V29KwbKznITzSM+dCrJ
5CCWRCl7eWMYpiVeCVt4/PVSZ9jv1tJas+hOR9wwJ3BPrbhgw0gQxH5sj60dKGD01yDJ1spF3tZi
yU20oESs4svbhCvjZ6FeOt9dDbLfYNwSMSl2W6ruBZP048rshl1T1va9YxQpeSKgmhiJpcStYms/
W4e8kM1e94CktKACBTpA4ySymsxW0yLpyjFEuagwsxn6b9Kw3jWvU5x6glyXL+tv5/QBZ035uTHV
L8lN0L5pptiUGGnpFtSwhnVAiFBjOZn0wxsq2ktAr0+/NDsr1WpBAVQ/P2023QIMR8sGjLEOoDIt
M9wQB/doakOYBJaRSUSVjPQzBptZK3wHQU7PqslRA18zYDj2ARqnruBSk5o2iyib6q9oW+aXTVRY
DufnO+pHA4slqawGmsO6Zs8o+oS9aIlS+6iNSS5BRUe9mdT2PI24hVpG79ZZHlCABXgiSfL4r+GQ
8qghCtFvq3ahFZSImYQN0s7SSZaZe4s963C/nR5UXPZnkgGI+MOi5zmvVRIGXxeErhYck8Oc0//M
NpobhtM37eyBRkdjP4wBac8Sd0qC4w1o0PmBKQM62CyhEM093n9AcxxayVOUJbpqEQx2YYflFQ8m
0FT8h5aICQpxFNsjt5CyxrCSCPqbu1tfRlYwmTk3te1vqjd01yCZUIiaeHMq9hou4cM0hxZFWeo5
fqZMCK1nvYcFMZimHtBBHoCRuVPqO1K621vMpvtAf8MfrBDd0cBohlEwbn8pAV2gEkK0F5bhBoUp
m5er4fgQh/RuXUS0vsKIoxzYoc2oJn6FhZuI6DsBDajTQOLZJFGd7tvQVxmjPJUqnqSncwOnImON
1ViJ7I/n1hZk6gi5ZRL67IMFI+5JRQYEpl/As64ZCDjfbgA11OMCSia5ldV48b9gkdT1R20m+7sd
xh073mLH7ZPR+1LmGl0wl8mGd2J5JQoASJRNPWlvyApIB4oUTMaD6t3JHRi2sMVsopco5i5LJ1i+
aKroI3ybbCJoT5MhECWg/Qxcu6xQS9+B4lLV/Q/losxLcYVJfpjHv9iQlK4wpNy4fjIxdIdamC2h
1t8XgHwEz1Dn5abiXboDByHUxuc2kPtOkU+d735P0OpqBgWN/qT2E1jCVWFyImLD8rdDUeo1lz/A
FrLumnjG7MYnroJJyG0LQqU9+h3bGMEY3JR3hrrVYWS7CkET1PM63+2o3a28mGF2ge205Gqj2gXk
3zuMpDdvkDMU3IbdW1Z2H6NPLx/0cFb3i1hRs3yG3l4WDNXOO3JupwZYeLpyd+tg5QEIaY/r9Ug0
3bSqQ+5C3gMFJF30mzbmeN0ov3Q/wcpQu3fbBvPA6MJ4u/wyKG9MLwo0sZQYt8wgHuysodwXl3Ff
u+rU7oZbLPjeXA48SMT9faCMQCYxhiWnuiVmd3cdtiEEeTbnU/wnC4cDLLCcn0gluOr9HEN0B0no
NPK+/d8pdkyTHfu5JPp1UTdrat1DgdmEXfqf4CQowKWX0jbG35AM4gZMParhr1z9excqlUNmY4Hq
Tnc5lPB2husVYohvekLjHMf+4njqHdgxFHO255lzO59s6o/uVS8AzM/um5pSyDZnmhxrC6cqfa1o
ypWYkPTNTqcXMpmmzqyK4qse+CYoPUBqNHJTfCnMIZJus+O2UfmCwES7kSifAr0n8z4n0w8+j6zT
NGRM1kPzPRUcVP3SphqSjDNMbsrzdiTxVUH7dNJCB4Rd1OVeI5udEJ3PcTZeVzCr31UyZ4s5rfbV
e7FL7hAbGk+TVjq1xYVROD7S/qZ5TqemGICDb+uM5TxkgJZT018/oPYu3gM6eK8xrGW+UfcrFm2B
zXt3Bh4MKOf57IvRZAUWJtXAQAwY6Ve9M4JAmNKUZTbGES8a0C0Om7thXOEaD3NC11fu2DH7tV/2
TDHchbIftlc757GC3SDlmHRti+3WkDLCwQNiStZK/ki3nh4blq9qndt0GyUS5IflNB2CvjDsIJEc
xVOD7O55qqsnZFXJl0whQiHHWHwuSZdsamJui+tUrNF2RevIQJGf/4ZtbGSPDWWGsRAuQuGSQjC4
2Ia0CXPcObg5FQq8JDXNkd7bcTCfngoRxoNzwdP0tZ7Jbab6k9VH//UA7sGbgzN4iayTtfub7R8O
c0DsaJCpy2duvzZI7Ar635iOjLNTsvyfjVVgb4xkhL8L1v9Jdq2Q2104XouP0srdi4WXxwPSb1Q/
Mrbv8og7sx5rhRqSV0fNk9dobEPlfI6mqpbcQVmXbtavk56TDMJi11WXn41QuUAlwL1KbKNKJMAE
LoaDTnTy3vQ/qQ9RtKVOd4I7UdPW160deFbNWI9/xkijRKvjAz/BRcCc+71G1cQLb12n663+H0Sd
44anHJ2DnARgO3bwpFpdKsOuqIsk8RklJ1yFZKJMrC+7Cs81LU+17soK1jWAw1tW3awhTpSi4xuK
bvrp1RJkFgpoOtjvTYLOoJNLROqEaJiv07Esm1OELLMScX6JlQylVpVjzh2y55l6dqn2WpQcoqas
kE9DxPliKdVThHPW7dmqFMzWRRf4VnIqdV/9hnE5+CCKiIv6/x4V4GU3LbwQ5LaIuXT+R02HDPN6
5DYu6I/ZQINTGvI1gXuQultfBqjiiL5fRdlkkqRbZjFAY7Awxrkww1REGQwQwRCwZ0I5K5QBMTwm
rluhCXu6mw0MT4X7/USx5qQUvlB/XHuMFWSf5HM4zkRAqYDPDxh660aeA5wM8kxJKsZSS05A9IyF
lpBBiBrTVQZCAGdB583dj96MKYKWipEuzSD7MYjs+LajBv83/H+RNvbc1lzyQz2Bdfo2ZfcG8yE+
ofUHLTqKKwUU5n3k5dlMcZBkNf0sLkaCpYogswGcY/t9a6AZ5ku/1RAiDo7F03cadBu6fzMC5tJT
dQTqeZXA8UQdH0bzs047DGlJh/2nbOxaLWNNoVCBKPsdB6ajsEFPrpfr96UqF6TN1SAzP8i6ZCjs
/qAVl8AD6dbt5HqA7rSoEKWHyHwzHKaarRtM6xVAsmC2ktiYrTU6mUdyrh55+ATAez+mcCtuQyXl
ms7AT8snnBdx/T7wL1Wn7qddWfA/42yawOxhozBsoNPRH/FIKs1BKPefAM8PJnPki4oDG0CRadpV
wEuwmgEev+tmYaO9mhJRIH1STzpbtY0avNUTe7Ab5nm8xyjvu855ie37d3TYxlUX7rAWOKyy9VDM
mEBFGFxMOArvPpgHdt8pLP+brQgSOLYeU43ai5MZTfI3vx6l8IVfjD4N8y8iRNqHE41IWFdSmfqo
JegimVfGJSA7b5GiWb9vtJkBDTRZCtL38NEr0tE/ql+ZulZSK7LCss5VtlahiJRgrjrT49WVTPqW
luQ5CxKgtNoSunp9oNWy4kCUr8dxORz3+x4221DHrpiry1pX1mFcXgrs430BCiAnGbXFk2sZjTsr
JdeWg1zLw5LTmtflv2uf2O8WSrGZESTjkPQ3A2Hrer7r7+XVs1SBIaYSPevIT/Wwwj3XblTBrkww
coddhpSJslWZCr5gEeVOirT8X6pVDoRewZhX7QF1YXzVGyPc0e/QYkRIb1t2FL6CJXrSubUP5/UW
vjnf3UwDrmovFn1NkfN0+HBJpnEUcQnAvm/PUhixHRjlThWU/21RbTcEFdiYnDKdXygsWXBfohgs
ASzOuBAE47mP20Xy6Q1k7RFjMJ4eRk0eNAUCs92enahFgd0e5iQAaIncQgryDw0L1/ChIOf20X36
PCI2NggYy89HF8pDqeUt99SQf1YTAr00FXhMs9sy1zpS/gIRnU/dEuozGNwy9At0RIlbfOUVPMUW
foiHazowbN2QUH+FUj2BBydSw4Ll34wZy/qVIO3WxywYTmCk3eh8XUbfDgP/0Rj7dZzuv7eYQcYH
1G3VwpqBmrSiechVnAYhUBvIOJDEW0N82O5JfRfKlhpexIH5qOehr9DGlkhcfssB/9tl5isJRWT+
bsbXXdMncC6N/59NUvo5KnrixLwchQrekY4ikfb/UlXUSIziyyR62BS+HL0GC71fBeqHutTiEcrT
CAk4YH8JzltuD721l/Bntv5SSo+UAqZ6HoLjZA3QCudKk91IM+LAZdF/VEcuwZto2hCQ0l+/ypHe
cmIspsHACUqNQyHsu7OLRM2bNpEOJYE6uDalCXr5ScYkfjS/+r2P10h/tGUD0SS8zvPaw1zDMojP
21nKAoYyW6lFGXde+u9MoVtuQchfr0x3ITQ5kx3w0vMK8GnrC45S19YbMW4rCTEExQFAAnNVvQw7
FWTywvh333LfMsLPSbBb/zszzwG+hY1VGRGTADNGT54Q+67DEICDNKwOaYVJKVgOmtUPnMSAhyn3
SpV5uIMJ6LE7D8RCzmqXLYpZZ2QhLFSX/bFNtu0QxpKA5h29FOS6yYL3L/ELKZj66lLYpC/5r3Qy
b1IJhedNJarlY/a4I6uE18Bdg5i3BFEChEDY3O3vR2GnecXys/s5WGiMH3r1ow34fDzw+RiMS9x2
1zPbJr5GiDGC7jbSJkwowolDJ2HJa0YFyhr4ZD7O1T/wjCUB8IfuaB09UUY2HSxJY6gB1CYKiGAP
nG25bHcbhpmFugG9QmtKqcr870PEiKPA97QJkOz3uAAF5q4AIoOvxKsKGFrnW7rw6OC55cetgvhu
aJRv4GbT7L3WjPzDDkSAfgeNzINPJl1l1dhhSAtJsJqA2cP35c4o9uNSTYwEy20xs3KftzQPVerO
iZtIPK39xNkkXPKV/WY09f1eMglX5FfXShBdFepIqwdDUafK4GFvbF0LOAkhr72+Nf5o+kO8mFnU
7b/KFJCpa5k5ok51tWkMgjP9pRWG5NT0onPQ/QBY8G8GdZ1MaRfjYG/hC2EtQ70XcxFOZMKDPhxy
AX/1AiiXLfgG++FrXApfQ5RU2012TS2DQU5kfT/fcKtAoNkOIem0IqpWKdxbQoDHx3K9icaayH16
qA7VjAhh/Z7In8DzzOXhyPxc9IZn8MgTif7TKBHaybn88fYngOVhEWL8LVo62MAA8mMkBuQHvl4d
dawRPJ/BRnYxjViIq+kDGdMnd2fDKbBVw2DvIv5iphljxRtnJhe8v98fXxl4kDkYvFGctqxQ0VnK
wnp/okYq9/TG83PhlFPmKtZHCB1NORedNxunZU8Jgj2Mj00jbShToX84Ili0gVNgMl+e8Z3/Fiwe
y+d8/3BAzzS3wcMxLxjmv1KIkgFmiN8ivg3EajYCV2WzxpzYJ9feaVCSKm1evX49k1CdQVbh8Hl6
UUZ1D0FePWKo0kxq1mwmpJgkOOOOQJok2xzKtOuV7bN4w3Lrle7DGWv/cjUPXK5Ye1zWs8TUwdYu
6HiNcC/01BFynKqw3KjkNjJt1s5VG0wG3FK1ozRuhAjkYhSOoSiRnhyASNOiVxwnkwMBhhMtjCal
2+udKm6MUgFtL79f/LsUsBdAUDlB/LVOWo/WtX5ScgS67sJvFEQr+3oo2Q30qSWilxuw+UCtssgq
8QGbdQ/Sa2V42j7b17pv+6925QGllQs0UoZBaky+UYV8CRjnYUTKO9bJQOPiF1A0xcaukIn1Rrtv
PWvqyqqIYixv5hmACb1WB3evJSY+XRWY8OYF5nxAdFelTaK82FjIekT1uIK92Xq3HN/+Zc5W2SZI
LXTEI0Y2G68vloqv5k/pMV3d6zs7YxOyAV0Yqshf06Vf7uzGJpXvJvsNrLtjVofRE5T3uc4W170L
5jt+rYt5rwi16/Pu2tIb7lOtpNff/nfW3tPTi9ac/ktMhD2iEuMHMtiWN0j/Be0A+ECWhfePySg6
qZiL6OeRQ0bJW23th0WbHL6niSHHGCj0E70Jdlpi5on9A10OCtTDCJdpqo4u4OE7LPuPVvb9qXSv
H8yKFitLoUOti+qRmFspe+K85ly9CA37w7bJZk8RWy4PkR2pcqDXCI/172Ua4XTOSZ1iAM/zMurh
wmNnM/tBF71OB+Kyf2FghSvB1P/Axh82N3gBYvr33hk40jTdxFml2Wp3ZlJao3SS+4byudm6L5E5
IbAaKoWVfvKiD56iDw2Cr7Zm13Dfc49PGgpPA/LO89Pmg3/N30cDUXx36o1m/u/HQfWJHCumtR4n
af00WVpSSqXNw1b6fMocKQhNVxqNI7qOM+qqLPPyVrrcW1lZS1Hcn9RuZPjy0wDF5gTT9WAPZX4r
GWALqGail0su1/uFjoBYdParxw7ESFhf2eB90jMpTsPOn2GJ0kPMA6Lht4HEcr89d3tgUR5/C5x3
oevGvEc9gDrWh2jmXZlsOtdIDNCd5VaqPFuByRj43or5SphxOM/tk7N5AjktFGvPR64tmaCslUCQ
ASQeED6zLmJgkVUJhRfQRkSlI4mYIHNT++RIAIXdJA5ZEHZ4A52CNVvjFw0F5j2aIvIDyMbBqzJ+
rXwkZbsX2CpYSQ7yKvK2EQB3c+RIPumZI4j4n7CbTk7ZwZCG97JL06Q7W/xwIcDbdYBkGslkTYrG
L8BM68zH89Qu5nQZ34lO9qcvt2Nd+6u/YJcAOpMI1f6ghSZhHQna0lqLRPX8jvFg8g0CICR+DpVB
RmkG/YxoavYkqPvcV9WlIq0c+8Nf5lddQWMueowjuDPJGrCx2Ls8rf83PtQ7/RF+TXFa1OUm/wfR
LlcS/0+xOWMgobzpcVqvJHW6BN2uknaZ8nnc0V1XkZCChtAFtFEYmwXwzN7VSrVEYytO+rMdn62J
Jyp4C+EkCZEjxSakZviJm+Pc+b6gZ1oeh1jyfeZBRwGB9Jh0f+eYq2Ic2qEk4UM8zU1OizfGeKN4
D0WJMOW2JADIE1DDopxHDzv316i2cBt7KVuFdJGpJgK9c1/Xjk0JokLbsNss9QiUnS0/yEgMcPmq
sEwdM4yuo2o0Czsl4foJPpTaoaqNx1ESWI3LinNBc2M4tKd87L7+LmMAuk5kDUTg6FcygIRULTAl
jZGs6HBY1VyhV2wpYzu0tPxyWo2wZTapZhokEWwFoVGZQNJ4ziiVfUqhLVEFiWm7DnAVfgdD4Vh0
apKPGNAVSfFD1JD/L8UUimm8iGMrsWaOiM6L5k2FAMfn/E5krZVD1aOeqwGyBmd7T/h6foA4dO61
Bxh+uTaL3/lsmBD/C1LEZp0SZMPYkEP15rjyxEHZPfKQBXs+WObYD1avYkJkbfE/KGFhZb1w/scz
B8aJeL/idQp3nfdmnnt/e/rzek+5KL5jtfMoyiA2evXebPolfo9uvRuSbtmEm6ImpBV7V8lafVNZ
6Y5gGsBXq5iE1UnA2n/F0GawqEdV8rf2eU8ZqDVKOBr0wkJB/W88EHBQlW9NXtOUxMAr7OLxMwRj
YylG//2+7SaHPjlRcLdjqjVvFIz31x3CuqgFGsbgDx6iM8dpXH5ZJggOpBTs56vPWhL1WD+TnUWc
zNLV/Vsa4dP1+batgz8aJxL/WMXtwEzu9Kqu93f0Y/hGSXVSi/BVMMDNKTAq/yOJ5rz3i6+Dq28f
lC5N5tDiI3a3uCnkmocxRVh8Tl12YsPcSXANqGTIh0lSWmkjLdU2u49gVWPTID7VjCiDKU13B8bu
YaEh9ZTu/uah0sesqt4DA6ELgFiMaUBjBX0RTgO32qj+R6GnJaLY9TtzJFnY5PKyx7gESLrOwDRa
4s9DTf8E7GxcIQnNoNLe5Dtg/WhrcvB+eEKtNwzPonb+E3kYpeRcFzjIRX3gmIuR8tj1KMfxNGpH
d42ZKS1VD1Ys4WVV9HuGQe8z4J6ZCCWtNP1ba336N1r0iQ+25vbz6IQKum4G9WZj6tAtA16XAf1X
sv8BzSxP0I8gNhlmp5uo+0cOefer1SAe+xHP79zCCNHn4M4vb+C0dN/43sHCeUp7yVHsf4GSoPpb
YQmVA5ZwCPw9MQCGPYjGVMTgkzJjGNsqDp7Z/UIHDA3vpCrB5yYlhx1C9/txIBTMIHDZNnWUVrdK
2Oe/hjPvgkzNEpceREs/FiSyrDboDsO0sWJDUzRx1wbH7y8EQz/U141Efd5lwhtnOX3sZp4DVk8/
j1KgcqBO1ltroV2FRb9J2gLt0PaRSb+xLvnGxd7mcvfBeNbQkISHjWmE+fCfU/4B0zCEbWmNt3JD
6FbrnRRyyt3aJjnYJ1aku7eANYxRcXbNkes0Bc8fC8eg6YfWXpxM5CZfbbyeOnQUilFtvPjH0JV9
VjpOw0hi4LPJoyn3UIG/OTwVPKdCrUP8oAHS945up4w6dKpdZSY4iM67KlmPt2LliZpEZW3dewGV
T5BRJ2dLeR54PdE8HZXI9pLZEaylk45ruNErm2bY9PuFe6G7VDM5rUDZRbGytbvxlXxiWgs98D0z
YO8wSYovIlQQkL1EO2nu4WN7l8EwijySi3ktwKzmxdlChGhAr8UCisC24wjEN6E3ISObxjPnShr4
//pc5eMoRFF4CvmbF9LzBKJs99NvXmjAQYGyS/WpNMQwlrG+7cF2j1ioTke3x+liHaDQuThqXxNv
ZdJocmMRG/eVcLSMPPa6TFEi5BJzzb+0Q8Bep2fBCEslEIq6zPTv3YgslnbJeadABHrulvlkP3jq
+2wztcNWS/MIX70usd0U5CPyN+dL4LH0cnV+qxg23iIq3BkGWYMIBiPVumvwgAV54aLhmBeXnDwT
uw6iRkMsh+kF+jEZAWBtsk9hwHTnhJG99/Xx8aiPkPCF4rCYTnp39gzLu3mVL06sSasN3zamZG3U
DLjoBKj+5YPDVvK3mMW/MyDeqhqU8dBg7NqyY8Vakx2kG421IC/giMe7wO6n10Xz0zM45om5eX01
CLiKkoC6lZMMbIWiGuIbnyKmCVBO7NeNkxIvQaWecZFwjdKIRhH8zrqwZHxw9PqtnXI8vzNwBAi0
OWXk7HGN/5CYLpXi1IPhyQ8fEMT+BpPofYBRJCezp6n6h5FBsL/aIhvkBD7/kEe1nQKzfeAbrGD+
Opm9N8JfbmxlIgUFueIGh06+jtBWsnNEwILG8z6VjjN/UeYIMCWzUjodOhnyszr79QLFrPxkm0aE
9CJkZgjfr07ldjErcSgOZTzGqplVD6x/q3aXRqZ6/o7TovtfB1ZWafj0u0jtaMxTwiyRQiOl8MB3
AlmLISZWu2T60ctgyokRcR64Obx9uy2VpgoLJDcHRLQLwsI2y53WNHFGeXb9ngfDCJFbLS72IsFF
VpXXYukGpCzjKNYbr3AL1UViqAhAFduRNJ1abFjhYjqAJW3JEX4MKKSdq4PCqwx47FyP2/j19bMA
Lj0fsn76eSm0i+Ou39G9+6/myrbPRQaOX1XQIUYIh9dGQY3HSe+NvcADzgmAafxZfA/FsDUPgSuk
gMWv0TWbD8mDKALixXZAPUELjVjrUks4AWvBGZVNUjqJprwfU577lpyVUaDUysu7yT8yglC2D/0E
fDQ4qmD/GwWLWGrUwNlwIdcefigfB3mwW4pgBUHhdKQx5YQhxgURy7zQLXsFbJEgiPQ0SXBhJGHo
9v9RqhNK15yEG/EjC7RUNWuZrHU6TrdWcCaXHq8aVoX+DE6avm0cw4/EtvgNA4ibC3bWRuv/Xgk1
M7QdEfsGaezFsA9fA8JF6IOAau8Vr5AOVQ1ylan5nPyfuAdreEReKvwrYxJZXrtkMXP93Xnhisn0
u2Y3d4xw7ChAvPWgDnpuJBpGVZ96nlbA49OhQqwmwoPlv/2873UXBYf0wVDw5umYeN2bHHiNwIs4
wa/9QyTWOUniSwlX5ia/9iouySq4fUEsrqGH5H4Dr9paGLPPh6WSE7QV3+QTOSCd/X4sBrHEHn2k
d5o/ZYNIxAkgQhSPf22sigzizPEGhBulMWn+GICGjApdT0ldjbDzQK6pyiNqR1RrWSX3Gemke/Ug
rQfMI+t8qvPzSSlBPxrxrn/RqRUg/PtZPYZGz341f91p1+I27+KRAWFcWxf5pa1ey1zxiS2keem9
wGJDPRbDZPvxA1mZxjHhwmYXxziZic6KXGWy3lldcuB5dGlyHUxtIyFVnnl+WHkWPrNKhBccQ22/
qZ2Xwh3As9GjFyleAeNaDB21tZEBX1tOQdOl7XC4meePcXAuuAoGieBnCs7ozAYqI0a1Q/YD2O4A
3AhjsjfPa4CmklEtlzd11bxGxJZ9kWxa+VEREI7IUez6lqWAb0A2xzNH3zgk/rGWeO6gXlVVERKM
VFlftsBhg7mlZC5XgdNbHd3W9XUYMVhlytDeuwgm1ptE/9ELolWtANBD6Rcbs7YTBxV29K7aTqzo
ga4fZ4WcSsZpSI3MwjzCW72PiDrLaTsTN1ozE8HTd+UH7g18abAywwaVy9+znOoNvfTnFOZcLPZr
fS3Yku3LproKoxRQp5pnqxo7gUjXdz47ITUitSgU1bb6gNzsnWzxcNqJdxPaAFanv4DY8M5bsf1Q
QGYmeXPlD8KN00RoeZUnS3ESBhyUkaeeptOuERAUMpr/yBb2icO3bP3F4eZ8lMVV5w4Xpug/LYN3
yGOSRAgW0gLMkRpka/qzTxD/IDKUDH3Nkb1H+gsvzxZg7jnAJRXvsnt1p9yLd8RgeMvRh0zrwWPv
/uvpIwoAnYSQ3OPUadzm5aUfd8DMEMZwzrfE66q1ShhJzPkjveWCf1WKA6ynsA0q+0NGgwpo+VQP
rUq+PP+TqWD2PdjLmIKOQnL8MRHH2oquskO9a7VXpYOiGU4v6Wz7uV+W+ZpdzFM4ThAMp6GZjPGl
X17YmlQfhM7H1VFvgeE7ZAXOiku2ubiVZQcR/Rj6VwVer7EZq0bcnjVWBAS46+phkj2MHhI86tNL
G3KEayJjRbTkkfKt92u6SEsrRBMvtLCZ0w9t15X/N68WuDyQehv5DN5J8mVMGIuCzxe0gX3KF9pv
DrXxz7H0FE7Ml5glXNyJ3r2aw1nTKpaxh4ROE9BRU9Q8qwRlIf5rND7z4dCFD3RZdU2fFUHsAPfM
mjLTmnXKa8cSn6HRT2GbjFuKQyUe71aLJhnCApM2C3CRRfREkeLsgQBFiiWWZJqkk5Revw8bQjMf
asd5hrNANl1UBpql+uoTY9TI1eac9oquWxbIat8d7CiLdg3LT7J8eLO0BNNVjYvKlDqWld4mvX2k
mtO2fv8XWtqiFi3/dAK2HZF6NYL/A54UWFf/5ANM4qqc4xeny59uNv6EiuyM+cpu5+SHK6vLPFPJ
nnpY1thsRmE1oXXVTroR+GFzll7GXP93E2ryxnziPS4Os5H+ZQJ0jCSL5skOzqQrhGEr9708pfDj
IUBKjeBjOq+/+dESq1DkgLInis3ClvLf1X1WIff/tYH3eRB3PqBrQCj9LgN+ChFoThhd5/cYiGu9
Ccr43ai79u71rSnGbeMbACM5ZkA+n8RhXNVfiMcsm3b2hNEsEuo2OshWDnQyTGGMaoN8lr5KlIt+
ns6faRKe54PaNqadSklkQKYRlCtThE7hEnCyHUJS35zVtAaewsPPgQ+yvSLJYvQ5ZPivXXrXdmtp
uO+a/61V7urvqOpvyvDbyNvI3DKQX7OZMbbU+qLGWlgzR39umvuIs5T4c9m7hdKboMpf+0YhJekL
gq5J+GFlax5/+PDu7bbfyy5MsVFKN5lShrQBTHVamRyCjpitzEWxSPv5iq7BgAe6OHnj1LyGMu3G
ePtv2F0/Gxt4wUICmXKNHKN76Gpj+4bD3Ak6T6aivCEPtzgdx6JSdwXu5XW6cyvuwKqZzpcg/1M3
Dw9kbKLrJhDe/JCIYHe8UFk7S0w+pQyZhdJ22Gvuu9n9aMs1SzoD43iBalJ8iNc1mT14LcfhjPky
D2Laqofy3bBB8uqoUcC8ItO88oK+M460sf6LMgbV+HKsOsY+hpLzaJPXzpvfmhrda6bFAex8XwAU
e9bSNKDcSMLyidXBYP6DzBKVOFrjjbwEZ9CbxFUREWdeeAwfMj7WsSkbUsZ8oQrrjxC8OCRzLzfE
3EUnKfrL0ve6bFFDWvb9UbZWQix4kewhwPMlbhYBfBbMZSxrIsVpMfQj++DgmULuPNdGM/M4/T56
eLblskXcEPEEL9+rX0+YSbIYkN0k+OZi79ruAb2pmbl72Eqx+bVkhqzlGCaubm/O15fjg7/BWYCy
y572kAgo2lPYa/j+sgaQlzEmwNQfYNuIyygCvKE/HNdj8aB5FtTgq+o7rAcPOiDx8dBlmOsA5RWW
8C0EIUU/3vSUMmqDrbnv2Fds+ISygswrIPBbdx/I8A3W8HZDEXM3/h+qBYIpmDivK91QhKC17S8J
x1YO7oq0S6v4n1GFE3mfxpFk0R0O4TMOY5sfUzEm76Bl7PdSqrUx+hwXGUcn1FGYGk8A7nh2j5qV
yAqbNkbOjZEo1PnrIsHNTz5m7OXm/ybweX6l1u6ZZSD5essDDyxQ3n7sadikI2OQoRLMgbRdbpTu
oHa+rT7i7NM8z2O1viE25yUyl8QkYNye03nAOKjwE0dAvwj7kREsiN4qrTr1j9d4ZRpQRXgrHFIZ
dBN0vaiqama3oZQbE+/o0bTxQKC1RdvTp0mJqS1ugJsjVypJyFHagbWTdqVar55nibP8yuvNZaAS
3FbQPfIXnnkTIzt3122/ZrmjdDnSrF/c7OouAPoYelVdxAoOLDn5RWjAzwm7SJwE12T26V0nTT3x
b9LVS0eb4UUQZO/9h8UXfopfsYKow48puQdoSpIDFSCfBwVJ11kjd0xh1qWT64mmD7OdhzTYoR8J
HhU2/3/Sdgsd5SCEIi+nddTuwcN6+lPXeJGlZx1TJ7mDkTlamDTh2ZxEcqCZ/PcSQuREIMTsbzYa
SHZB5csB66o/80r0DULrz7Xewa5neVBdnAhNtp+iXQZM8uHCwpIaOZqI35ZosF3Fj6k/Ve7FqBxV
FunIDYaQqCDEGPKgz/VelLEfbU916kRx3XL1O9oc+pPlXXHCBK7JHzgsYNCMF7PCsphMGeWVnaSI
qiKw6gOwo3uyWfZhiGByXp6gsFVROfZVjl6UIRwyKItB/dIWHdHRqkDsMWV5QuTzsc/xnL9lhlT2
7BvnSSFBRuTk7RLrc8gxFxSBbcRWXwf5rjwGGKBmNyWihF6zFsC0HRyQ9ZuV+GKYZ1wwEnNC4M+l
Rf4bVDZ5yIDSJMCsFDx0fiXbcP1cd920bc0S7PxWSudbqUvOYaRi+VhSydig12h/SDHOng1I8pZ5
I/wJdv3K4gGxVN9UhB9i571ZfQ8TD1FwmlvXwwMgmZSh9q7CDBmve8MJvuGZ8NY2jFb8Xgt0THeS
F3VkL+mfboCZxTh6Gz1PMUR/QRkiMiu8n2kzE5SYkqErQWvLs6Vj9wNwDwSPmxEQm/BAu+4ac+uW
5Zcex343X5lYOWQmoyc3oMkdgHDcojBpZHdtMmYP8Dm0If7907D5L3I+56t68gi8gJKHHwfDVJ3x
L3m0GtbcqQU/SPZV571jnrP3vRkR8VedryxmHW0xBg+3oqg9A9LeC2umcJo9t/LTm8uJe+QexQLG
E4yqkWAEDa+6ZVLScoFCY44DbLIgVMD9jIIVvW3KIxst9O856xs7qFiDulOvL+mZ9M+2vq+bcxyg
BuUWdbCf3SpJqXtF792kA2uGqg8WB1/b4tyA5oDdq4ENmGwgTxlHEDmRRUinkd4/UhR0+6Moteo5
6lG/PX4sP7wsJ5dqgOLEtxq227DkHUwq44USahJG6bDsh22NA4ZoXCrRsMDvkmmxm6fJ1dhkStjo
J8OCxo6KMuhsBF/F7jZmHJS2U75NSaAkL8N8/jkIpIN4H6cTrpttMpg/yvKe2WP69tjONOpmX6df
zfzsQjn5KbVdspDzJ1iw2/ls9rr6St6+yZrcsoj1BWNZXu/yGGwuyt8TZPdefSd/WMPb8wzW8zxZ
cxHefssWXCDujlInOP4FsWEZp245gqTW3hGfs9DhXu6gbYxlK0qhnT0IFwlq+aTj4oeBMp4kWaTX
b9vUcqKIEDC53YXfYm43eRPuoOTJYc8OPtOJBwP+FfC3vnNBQHr1elkiPl+c9wSc9RjCWL1wLtCy
QjAv3ok4JD3sbwpFYiTore3TSG8Qfmfc5BEQSgDJktfuykquJXIIwb4WwjlH2gA6C6D8jAozgvVY
j5WvqoeQ0JC46xzX/ej2nfdZf6uQKNKLdNexxIqWVeYzkHCFUzekeZxkf9dVzD3SmRGsafBUgRMj
74ewk5WWsas/No14xM3PLEKIc6jFnm3XvIzTc4g9QHQuV40BTB9WFZWyietfSWTFH2uvMldY5kam
sihc+IcuSAg0bVvois/65K225exwPTk4zDNa/FTv70lq2kYD9aLipQb9jWal/DgkaYapG7z7uJQu
hx7hBNnhBJcnPOWQI+iCu97OEQmKensQssmMY3Rr7zAk8177DnnGzolIVtD69juvZBKl+pcP1bl/
iOBtek2zr9OJ0kUA1OiW3VsStIYMcO+V4KS976GYVZ740K1NqHLTmzFrP0h0ybanZeycyAV+rXHE
dHXpDvpRwU84UtGr4ucKmjoK05VT0ZvnxPCa6DO3GwwR/AmhEc7XnbzNL7uBC0PciEtKLcRBNqFh
CYSy3HExrHrxmIzJmXnEUtpckq2CPqgl1AmgKbzza3ydBvnlnQmEy9qqsS/lxrPI+uCSaswN7Cu3
wJvZ+B0FT514Bx8uaZbu2FPUijuRO59rCeKBh0eksxuA4OIDXheiqdVG0JEGferGqkRIYIPqaYRx
NoWSp+ELaQ/uvytTKa/GFPl0DmH3X0V80smeaVpll2dRo20X5tLCoxV1kOHnCGcMtuTDTQfeHE8F
yLEgfpvnFupVJrNuLngj32m32keRJdKHO1J17zbGrdvu58Z+C3//QmXV985x/Y3v8CLzYhfr6Nb2
jJzjsaNEF4HjUMwrpchZUhzG6PsZWOT5Xcnnfmd3ypLfLZ4l2991hLMzsHT7CaZeBcttEEe7ySgu
YMm7sK7QZFAcqvH23aUl1nt5vp/ymoSCJlD0gKS77kP5iHhBpKEvDaVdrkLoXhxIFfVWS3Fn8v6R
kvtsBRnSxERWV88YKhLyPOOwGf/H4VKTXk2pjSANwTQ4xumXMbbjLfyvSTnfaepvVlrVXxsbd8wW
stcJdh3i/8Em5umOmr4HY7n2qNhZ+7PYnIfmUh10Htx0hLQ7Mdkzd6R5D+ZBHXPnsNN/epQD68Qu
V1GGdWMKTVmt+Zijk8aEORGgAiktBJgUTndxz6TuK8JWq/OQVUsMa+CA4OrWyyOrJzv90ubYXTYh
XYaKuheGHvBfeHYGlECvZS8md6ZgX/R9SKbjQIapwz7zpcBx2WAUCPLHI8luaKobnlsHlXjAkI1D
Mg9FpoeKqfRxNsuKNXdSi9EdXhsmV36OJz2yabGr95O7YgOLJpUGUl4HsSDxUmb+ezoDR7wd8HeE
scgcd3tRLWOU5Thw5cewMJgJQBmbbdrGz7szN5oT7a4F2O1qC1cP5jeZnznSEJika+uqHeBMcvH3
l0nHOoobs8HvOtll0LCBZx/bvfQF4EHuJ5vC6cH+D1Os+bjLHd9vW/GqR9rMgUM5zGbXokqApyvv
u+1nSLSymsJvWBRUqREVzQ1jo39QJDIkPS7dfwWFOzDdOl1RR8BSjKwexx3lDrBsrMJckEYg67G0
aFwEt9+zgr0cfqZs/xP50lESzK1eLu4f+Z397eFeOwD7sjE7vYckuFz7nEPutbgmv5Iw4irAwUqn
GoFPPRf6keAsfwWxT78FlhyHjQS+DuUjOmtL2bfib6VkeAlAZuOJcf85hxEyatAYQ/61afNIa3GI
LE81zD+72WNFn9StiyPWzY65qbFhj3nwws+UQM3qzFfXqyuKscAHwrWxcSZk2WExxUFdE86aYKR8
0f4RUIVmbx4sGcxfi8FWS15lj1yohA4jg9ni9yZ+xtSPN5AOTLcx0HYDCgzLeqCYFjpCJJOTyL89
Qgu2y1K2dPZf7uiBzLiu3wQbJAmxY9uziC0exVleQUJQcytFvvVOGa6eNFozjTMI+OZIk3PsQ1n+
aQ/uNBVEbWaNLRwvv7O82iKXkYRljRElSYYFIOTAMDzfsv2g7PyZD5F1PfpK0hdLRNOcdGDGCXQV
7fp04YBCJPqwTPnLRtZaC6KdI8HW+74N5FJH6ASVSdaVbTMEc6aRguUgefVqu86ZJ3ChBAg/4FGF
XUkkm1EBReGYUKtyPEtl2kpRPDFAwCFvdOlM5adtlR6nnIWM3Ytdv1giLRWnUuIiC0QA5k2yo6ki
O4YAbok9zKLutOwMEN3oWpyd9uzWkPmpj0g6JhSl/O1ef2TCpwJMvBHii+FxSnM9lpoW6fPKOqdh
upYpuiCqBWy/+G6Eg2ESY7PYE2FA02i6LdzxEr6Wu17M4TMVb5/RRmVmLW4mwBF1f5ImoZsuKr6p
ykz32k/GiHXw7oaVDbeXVwomnx6ENmk4dGRKWIWbC55z34TJJyl59CQKiIsY2v9zLTuMsRFSmIAb
KF58H49l+Ul7Op6SkkcEflj0HN6GCO3LvK5RIimR+l8wQrIRZ2TZya20/TEC0Iqt3KkzXLxHKG0U
S5JR7ql4fTxaU/c97I27bREPnm+W+363LDIhBpZnvZP26jjqb0vRsQjNOpglZbR990zhwQ+hPnjC
u2nIHOUIjKawd0t5Vl0XfaL6t522cnnphPjWHj449QZVDwFue4/kKFDkgCz8lJ+rRJVxJcquy2Rf
ZjQl1rUksUaJHwloTvC5AWu1YzJjZSFKhxPvpjudB0uL+/dMJB74xyWiNwKFbKmQdDmJ9zcZszuj
dccSvtuDFuI0RQh2R7rxuReAYzFzBTOtVN53w0/OnBsQBZZlbtUwRbiQbCOWYkjSTza8yRgm0GJ/
NQ69xp4cxglZJpX1KV96ddxW/PEIxqSogp0ACeeDiivUs96H61N2DQiERWuoFjlOzXEMQvfPGiNW
zXcpqy3b5KGM4nxQmB5pP+2Bs2WsIwoPlOA6SKYrMt9VNBsb1ogKUxhPBjOqERi1C9Fe0eRl38jx
hXWJVsH+8No6+x2t1LW2ezlKTiZZuiTjGxMWxS5dSbWtRyJH9ttl4FkZT6kFjB3/yQFNYCMKBFev
WJVcfJ14Mmbd+If+56bgUA9P98eeOc1sFCJwk99Ft0AX4sa1J3E2/weUArs1y8rnBtiJCBhh1uiw
oI2BjXT0ZeVTLfkRfW3Hs6Yhx4vEZKg+UeMJXWoE7a3InXcVVyCCntKG3SA1D8+nxvzLvExyGqQo
G/Zg/z8Pht6fofcvdS1vrEPGxAryexpFxbrEBTxkQZi8aJ5CSwO4WyEQyrNacTS3uQt/zvQ4eFkp
0MxMMB4OlWRiVUVC7/ODnVFo8Cbx4v142sw77alH42vfOwiY0adMYqVhOSo0fMy/+StVlSm8G4qJ
aUW80gT9d5cRCzlWC6YgbIOJS0G3+IQvSH7xtOA0mQFs9oZ2Nwqk2p7NGSqlj7cV5DzrqDwY6qKb
zVylIzhSUigetG4jE/emWvWwo+oWvljYrrtFzFCl0tml8H411JBS51A9p6gehpGxn80LxFj12ohm
DmySkrFmr3aihgEKgvdcKtiBLrfkl8NH3cgLhO7LwBUK0xDr+/AYYydgLiEbHxaq8C/NBJukuMme
YwZRD3ru5Vmy+fjxIN5jsc/68U8uoNoOHr4auYzsrKgHgKleWjJLkA5fd/S10VV6lBqWchtuf7Jl
CHOZMMiOX+cQSqjocnEcfT+ZyHvrR3/6KZ8jseUmehREMn4DycoTxgKeqBLoy82Pr5EIldP1J91B
KlTZw8VblLOqaGGVn4DAw/F7Kc5HKMrpSk0jX9QW//U1uic915Uisi+2gR4vFi0uqn360Nkx1TMz
wrQ2P9zNzvl5SXLOZ8cQCNhWewv0S5vNNk4a86e5cbK3/6MUPTIbTSHexknDNMe5M25wkEz+NFGz
YOWMd4r7mOnwksqQFxIwZT81ptjjrpB1JDJArWsKXhHNkO88GnJETi8msDTJAHm/CJp5qEdxrAvz
x4kB8GGS8JjNkFpKtXLbstb5f94iTNbcfTceogUp8cNSNL0FDZA4gQkPG52XGQF5R66CSOdHvxSK
LZruBb/EH8tHaAOZmvKXs5YkQ1SzmscC8rB67oGSJouni/OiGDoW6kAGmWtOJUhnWmbmCOiRp5LB
6Kiz47tiwA0JMFMz7yP8VBesQBUMGAJKhz7miLWWF+PYaikMytuVwNHkaVjwLrBdETm6a15LxELq
4PoWvEmH6ENWIMRq+pG/R6Q1/OGncGVzbvX+e+oQoDV8+zcIV5ZsSCUQD2rQk10HCmJCGF9iQwlm
mRrqQ/V9lio1SzEVVBbSG3KyVN7Vtdj5mlmb/ApdGXIkcp7quVo8gwH/3gG5WfGWTVHBrCpDkEH9
Ku+LeXiXjfBI9tyJgYXdSshkdAQPVO0++8erLFsL3w9oif+ROPLgBLWD2sMbO191lMsry6Tqr859
n6DTcfFwlk69O/pPONktDJ7zVl794f+iU7k/b041ttzY9C3P7Vot8ae7E1wo24ow+9U45w1X1Rzq
cUm16adKIzg2Qt5euZbB4QQx0Zk1u8DeFny3ve72UN8uW4ppiLBo8p71wmD/E8dv0jus8/j++6Fz
xllmdupSEHV787KNBO7fNVijwb/+7WGx8nh6BXRhpHuqZ2eBbFv6Q8ofnsienuH31viulGeDXFid
bwLBOmdoSbmMc2GMxxOD0fLN7w/hJ066zqiYeauLeqlKGKFatvv79VlFlT7K4bTAs2pdWwo9/2KR
L57bfeJYj8QyUxuXP6rpmxhN2mKxtsf8I7iCvx29V0MQ3ryPMFgx7+X5znRFr75Ow4oRR8dnkvnT
9QUasGZss5uxRxSSxKhrnjutLBG/FP4hXMTRkHmEpXtKt/4tZhj5yLU0Sj8+f8I22ENH5MA9G5y2
m5T2zzWx0r8v85v9+A7EwsHASCr0zbWgBwfjfTOZxurc4DTv3ucrBYC6YhEhVkFLg9yKO1FrqEn9
6dCG2f3TV+qXDEb4kyuMCp/i4p4fzgMZX+j7HV9uKxf3352v2cxR3ctjc/N9aEu9yOSzxskqij/3
lfQfA+vFOUue4v+tDzDIHakswEF83/ODxHC6+zG14iOSr+J89OL0OLc4Z+9/GVYL2TaR4m/qtcML
o5vFz9sW+LyzBQRdMutBwT+Csq0WO1Kt92tvErqX1NcRnnvFQak3GGpmB9MbgHAri9nIlFQgVUem
0DtTR6ev56Xg7CQsEavSJNQnGlTIjEIP+8TRTZjuIW+2THWak6vSqVJ/+rqDky37H9HDRiFeYGPd
DdijGJe+zKVvlbqOa8SPV0NwYmCa8mP7jueLotk94oSpJNfXt+24lsqGdE1aWPK8wGXv/T5DLOWA
1KdCD3iwVcLqKQFwundfMZKN8wsmT8UnOZk+xKCLylf8QlgyMuFGQgOGAdyfRgJgLaZ+29B3Wgtb
tXOmy+lRNuEvtzXysiA291U94+UgkwqPxrgfK3u4GrshbgJIYdp4zXL9RG7s5ABWjOC60XJrv9Ez
sr7Og14aOmp1i0Uoa3o9K3NLWxfd00/j01WTALqYqn0mO8IVmSD8RTd1N0Ph8v7rQX+2auoaPEcd
/IhgXkezKc3OdEscHn2PqUJjzK3F/ADyN4tC9WikBcHMbvB+N/WuUnGO6vbqchFxygHpUrzwoRIf
4zJkrsCpIab4pIEVdOUhV4ioWzgEWvedYmoD/6TND0x0z/w8DM+gONQcFhjkkxXyaZM/JalTfFfL
bIDLLwnQ7JfQ8gQmvAfm7sDrs99Tg8DLLngcg+MZOgofq1SrV7nRg+Sh1WkDqAfck2mMbADj4VVI
H0aDphDLuRQhFp28DYvmBkb0SiQwiNVX3yOPMSK8exJ1Xn3BfoJPYaGUE0qltL5heMsxDjRmBqFb
hXQvKr6QXxQ9EjnaNOYREYmoDE3AV5tBzPzIJPAaPnab5OFM47alrVaoveRxLUbMh2pnZfsk/cMY
E9COM1VVXyYtq/lBlVwY+ODAEYSG/fZPJTWZBCVT7GaDf398j9XzcoVpmy6fkTJ9Rw9/egg2MDm6
ndbVLI2BWT9pafXqnswVPqtjVPXkgZy6C3xZ7ZD0XmJ9FgR3U8Rmu7LYSYY6Al3bvIFeN6gwEQUQ
hjhbSyK7Py3jhWswG2Cf0Vef5vzrzDEhoUNCsKXpk5lx9yneRwT7Yqv6WVrZ1H/esAuBv4bjxbfE
h/TxX6eQ/cWHQtuI/FQq5WccDEYGj2CMA88aRysVuYzHSvbpyv57JkBUIYRZCSeJ+uVOBItP1hBo
eeGKoF4m05jo0D5aEHQZtynV66RAdJ1rUyT6R321ToT2Ler1/TBBOottU/hnQqK1/fmpEXurHxzQ
26my/jeOuOSjU57xNjYPyXZ3+IsSWn1FlwjjHD8Cw4r4/zsE4bMmTW/rR8445j8jPRK9/lI/n7/2
LVv+7Ng1GaQfC5gjPQZl/v8b3RBhgtaNrZ5xFJb0pDrhyEgngvRoCfsRvbimZklNAj6dFygDTndX
PmLqSGzEDbocXCgP2ATciig+g5scuBhItv9qBTS03t7z075Nx9tIVl0n+y8A+7QzhenmSMjTacYc
S6P9oBSFpFo6jBMLa8fp2zu/nlh5szmUa2bEU2BDRsaIif77EjkejXu3pDPVdnjLdwb6LZVYCqb/
t1ooNVnqlNvCjRngwcdD43ewYnwA9bxZ21QgFXteYrbZmRb4D9RrmODb7aslXkFCFAQV0ZfMsDRW
sVlf0R13XF5fnwZdzlzuNInGRSr11ccZrnHOSYn7CdRnGX9vkER8+Ff+FX2d1+uwAqQI+GnZ8VF/
8U63aO7nk38XDP5QCk+WmoiN7RoZcbvjAAtv8juelfxYS0FTJal5btAuDuwxoclTNkf2dbe3GuKl
v5XuVD/cIZ6hkXS/F6cTJyabUJtGRp5kgiqecwMJrmNrNVA/z3DJraVIqbn+gxSFFQUW2ZPhQOcZ
EeDJ83rRxf6HpouUfFwmB7N/tzqrAxIW/qBWWGI/czduCOf4+IG70suKsh6+56w5Bgcn11r1UuU7
t4XM+Cy9m1jMR/Ds0x2A3bqMXsaKn7C1v79/jfquADIYh0Ep0ugi7vYFarJZbiiwE8epS1CRc80N
5y0U7wVWgc6W+UocpULL4IC8+vF5uHiWwv+CsmM5lDo6b9N2oEG7XJV6VYg40ZG40DQ+/3YQtU4Y
bYqmKrejGpCRTMBUfVvilwLdUHxC9C9L07yvDmpFuxP0DnESB/qa8Yh/SwsDZUYE0nsQmuvz7jTV
7RFgGKX6HN6xEKm4qotykOwk1iJx4lFnJugOgizPFyMNtxCMtkWiriIoj/esEiM+x/TKPV/nK5Ie
SdnMvYm7anNE6YxWGUXRODu3HSYZlGFgTMzP6M77n62BUQ/KnwQ4q4fgCuYSj4ydJTMxtYWg1cJS
NKrmrgXSf4G4JvF53rN1w9MAIGK3BHDREmm9Ns+ENhHaFHPdA79m988Kce4xUWzIS/iX9T0URGEi
cG/HqVBCe0Ysq2ZDwJ6n0OacNgPsirZD/6624p5oXNnAUE6YbvJrhcnACAfE8HIO5Nim1bX0449M
bL7WEc2bmzEEseLw41oc68283OZVWDTmWAgb+KuXVBn2RaPqpmitkqoNgf5SztritnUEJ7N+/0D4
pU0R7aZgiz7TwWa2eJZ7+HVD8rg1y34ACKJvrXwe1+8D+GK9m2I54nLTIXMUWm/8N5ezCvpSjrXL
M3CKw1EXV5MXV4DAE5YS/K/sp5iRVw9y5vUxtzAMwOuv2x3HobTFWQBriskvSqP146I8FHetBSWm
nCFNXzGDT31FLcN9/RqCC0VkTAQQwubD9uaxHsxXctSf80xJwG+/jCqSbWn6MEsi1Gq/ITBIAfYj
YI7G49TEcEjNdvkbaqH1cKvLfMml6wR0RylqCnewYVG9P/0t9+KhKw5rLZiqybvZSB1x2PgqS47b
0OVKUXlKy9KipueLraqTaMiJJvUpcSNBv1BeSK0dbPTWR8B1ZqN2tTVZ4BGC38ef61RLxzaNkUjg
y2JO6/kcrMA8h/PbeKr35BDZ32nXNQFd1KEgmaD6FVJkHuUTAVU4o1bUAhenqFkU71TTtQ5SLO5R
9Rx45pvS4zf4yt8PPQeTIHx5FAg1j6/XR+2tZq3SG9XauXri/knQKPSI9TUIBdV/BlFnPX/diuyu
WqLp1A6amQQpF08z1cH8ouFehw2V+qEQ+KC2GaCheLRmLe6yO922zC8D8k/ne7r2EmVt8fRkJKVM
F6K1Gij2Lyk7FGWKaKH+js4ecXpAnHmOAriq8itl0W2FYBZELRN7AmQTNXUMgiL7+w+/edmUXUYY
1bL2q8lf76c7X3efjMe18U6WuGaZy2VkSYOa4cijkokvJKG+fKLoYLVUbQuI4M6qOvU1SWDiZay2
i5wk37UsM/X2KMfsR5wQKwRrGplgPbWhj5PLHbzk01XTBxJA0F4Hj7e6I3dxdf/mvNEl+8sbUSQh
6LOt4EdZ9IWzFfPLd99SwN2tGBoDx+xyGoR97hr9dj6b9gvxFPQZIUuM2+IX0oa5m6mtb8N7WvZj
VMtrpCJTRVKZIxWVOFKHfOq6CnSXvqseLMGBi+aoNLEAYT9zzlZIXqeK6xBH7mhjgcaHaep3RmEi
c+9EysLw2Xj/c9vVySGXGo/pjF4UzegyzQgdpZLfsF1WTEKcZph+i4Dag2td569aYCCSLAZh9uDB
2KTGaHRNtUb4xU0v4aJT8Gsbmfg0xVbVVZD9r/H+qH2QHBoirkNKfm56q6lowq2S0hn+ZSE8e29t
9J2yu4B657Z8FbhxzRXZrTWNOm0rvU51Tsz/EVBb0yxBb0qDyr+jmFC+oalApLUn7lnWJLMTFmav
ZTzrPOXGRiffLZN2W1tplbTNn9Rw+ZRJEhdt7ksgc43Yc7BOI0Qj//Y9i9SGwEb6fTwpvcCqjt+G
zPErqto5Crim4UHRgfeKQW9uzelJ58fjZ241fwILULaC1tBMkiIhiftt3iKgyTN1eFpkVlb/R0tE
S7DPhpGjVd8awUNqmHC+obVQhUzCoRpd1szVDhPK+0GMpRa7V5HUckZN9OtrxXsaTZVuO6PwNIkN
VJ+wufhkU6HDyOcyOzYJQzhfvyE9xNR6TJ77QunwMr6UvFyP3fO7OrWTtc98Uj85lgMm/qPnGJjN
e7ON2XZND+z6IRT6nXDAVrtS5WGWzoTaUkqKjZN4jMJ2HrldR6PLKRJAHmOyH278zkGTOa8EXtr6
lmfYkNLvdL6dAsgJagGN/l+khlmixW4LrwaSyB6NJR7W0yLKm7y1CL2sK0t6h8dOjXdjwshVrios
NVa/rv6xRu53z4F+OBya3kDMK02TdGDfEJvJNOS17gulrYps0KvJ75e6WCVc0DjnCcIAUt/j5Dep
z1RHO+yRQv9ueivvWvZ/xvPgnUBxZwRx4JcSNnDPGyiRr7X/O7yy3TL/okEQ2hEL4XcJmWnRyfvP
7MRNPl8i/lAPsNsb6xG7X8gV5AwHBIwhRKuQK5JxdkaKCyp9lLDH6rj6WUglNkN2GMBkwqO4ysOc
oktKRdVLDBTP7Z0MmmWBH2bUMdI33PfigcJh3hvCiJuKE94Y23bCtbokqTCR1wxhwvfaLvUTbzGO
bNBPRGUUwRvlmYLlZXmIDx89tg6SBIqTHuf3gHnlNw37rPeAuyVcDo9WifPo7Rkoi7E8eSTumqqS
R6JfBxogweloZ3LguHQjd9CR1Ag9rad7UtHNIxrGjfhsYSw+jIALxNtSyJZqI7I4SUTtOiQTiiIb
lX66hcwgsA1kuvSsW6E28SkXvbbCIWMRiHQ4Qe3yhCVYMfGeiMFcmTelS8LPCiLlfONQpg50mBet
hIR09SEIWI4umpkZNJIGyC/Mo3ChXP5GmddCC6QJveardm/Tp/VMsDxn3rS7QQ95B6IeyBN4bl1l
Bn/05LKU+L4DMMJjOMTMQOV2i/AyBsoR1ye94xxikn1PBaFxvnVUDvUrMDT1RSq2s9A/zGIVjd3s
41WpNxqjNQLnAukAuHpWjQIcCKvezpHS25uXckkk6M6cysFxwHy+Rw12ehE/xatlqLGdnnVL3ZXc
jbLdzdX/euTRqAeX5QI5DEqZt0IbJ+zXGHbnd9F6YLRxyCAjtEV+4rqK0AHXAVwS5H0Z258tiT1x
9Tq+QxbBoJmS00I1cY9MGOT1e90O9II5HDG2w+bUlhbHiG9WgIBpsQxXr2nW8BQc6CPwhV6RQfKn
9x4eoB//nfQRnKYaQrgUQ9c/nFEGhF1MAfgEux/q81QFgimxBgX8KpYJbii3Rqfv0cGYoywaooMQ
e3Y4YaSDbc7zvDIkvpIi/tenl53p32UnjQKvo+Cqjix3IpRhSpTirpXN5zL/FO3YbyVd+gGllXba
bkD6MNjRWrztak9iwu0kuK7JnPuhKVtCM10d7CmhS1sM5hwEIAlzzmgDN86MQCJJahCFAbuoNvQk
w16Q1oSyqI9a4rH+UwTwR7Bf/X9XYe7HnGoVyh+T5XSRsWxn3B+zrGvcqdDv/bsHBwkfZtl0BGiQ
fkPVDHbjEji5fVjMHh79sN+PM2rYpSET8Zwd8yoCfdilDTFcWqv6m5jP+TAyY7smVmZX3d1wpxLw
Q6h5z/gE28uRM6vDZjqzJfJpcC2s9DkVQIcW80g8mMQ/hANnYhrpoLZCv/4HImAaP6puVNKeetI/
hUJRYjbczqNRWIlX5F0KJYDtYpWiixZkrJeCYSTaWvFvvj2ayGlzbDzOebwaIw7YNUu0CtvmpaMp
hmbROt6S+m3gpXMhdFy+8ZMeEwRg5li22e4gWZDS9MUoopR95vVftpb96IZynmXOVtB84q0P0WIG
WVvcRfCWqS4yogd3GhXHWeX2O2E0h0jahWE06q2uiucy4gtHTijzhKk8TIgA/qEiH93BBFk2jIu+
4jU5ft1WM82Ru+i3ROvm+zqB3u4O4wx3rViMYJhU+Tp9TN8xpfiYmtZaVuOS7lBNm5k+17K41APz
YX9eCprV+7aFugprgXppoV3C8ClWNX8ncQkHK+wSHf5P4cMXNj851jE/aLbmnx7Zo2Qj69cCaD+H
BfVggXFfLBZhwBMJkLpZ7O4bu3TwIusHynboorx5L/KxAdMinTYWnjBCmRQ1/c+T3Sr4SMSSAxHQ
90oVdXB7cionB//qItqpJVSPHbzEnSN4Kx1n24/i37WnFU2XilXPaBGxiqNF/jrcRxlcu1VMVo8Y
VmrlKS2AbSABqOhUQYDBP/piZeK2WkHYDjxmI9Vp694peYl9jZLxkMBJAlm0Oz5GAIoT9D5VJulj
50kCjjPfDnvxQNLNAKcDg05g3kGGwaM9ce27JC0Osq4Zt8N/L/Rw18/37rbAK+sxWBJas167bTf7
YJzKBUP1tqK8kIo/YVJ7bazqFjDTWU0by8REpbJ0bqluRov9WQ5qOGHgjxwFyxh95MPnP+AssxU0
dgWeBhNULKhH3Bilm8dhNhyN7+L/nKnVngnYdlNgZBD1m7UkCcM8aeXoG3WwrENLIvOhdLMf3NK6
gW8EDajh8Oruan99HGk0MzWJI9UBf2eiI0ntfvgl0zuOjvKWEWw2Onqcyazl6eieYFxx5qENYqRS
tZzaIXuqlg+i+acoEeVNIcxnd/4k/7Bm9CRcKu+O8FodmnAXiP/zSD12QEKbl2gmNiXZbTgQBeK6
WLFtpTTpKmZZ0sJGSfTTVfwPRipVt1knEpCkMAFbuusg+vwI6zOFLqlYx/R1oQMfmxpKsms40Fvh
KJ2igfWSrcZvBiMIiVKEozPPl+W7obPJOf0XD9y6NP8YMkdh4dq+ZmeDthXmYIg4/T4ppAeznJkq
LV06W8m+tfeCrKyrF7j9p/MjtZ6HM80ooUT3si9NJiq3+FaxK4iTQVBaXEsVF3QfjPHAdG6Z3plQ
SLOrm5PGKfnP0F6seGaWKJKgOt3J2b4iQvbHH41lMKX9s8p2dOujsYPWrsHlgupTuyqZK4zxQh8O
Q3sAd3vsV93VTdZM36Z1dyE6T6RLs2JCG2eF/Zg7qwdy1fed5RULcUu+l05NLixzOv5HaKiOVuJV
u0dJBlYm18prDyjfvhf5ajcB+7Glshz4aXBxXt/OlwXJfx/ojaIOayHMPxwVgsn7arpsXOlHXA4g
YdwwL5PHybYb9X3oD9HGlroZzfkjJgFHxom7SIVVa4cFOwsaM3iTEOPcYJWKdOa6r0XaAaST7MuW
BmKKLOs3wuUN8U4NN1Cqkyq+S94DA3Uvkcven+udFwJwxn4IebHoe0EjMpJHAbHxf2hkobDsVhQV
Rf8inJpOWc297+3hPMNZTTstN7L0kf+IbwE0kXY5lo6aCPEf4Y/VwKW1NiNuElWVGUTCu2GWSM6S
SjHKhvzr4LJccAwOxS/YMh76TXgHujjqnzqomc+SPAVz4rGwA5/fGPiHv0Zu5aPgT8CWuQrcZPbz
EV8oiGWGsZzJXTdfajqJMW7TINOzIiUcvMcj1H7t6teVR2uoHoSsdIZPIxfKN2Q5IY66OvBNGMqi
h0gDyKRu6nc5m027MrpsEyRCxNrmZB72V5nFT/PLecKPomjYSnH5skgzDVpzsMny3lyoPiq8U39J
iOJKgdR27hWENGqGQZOZh/iXgPyhWWFS7yXteUPS+NVP7gubno2Palx6dksTMCz9H7ReizBUO3dL
01220zw3j3ueRtVns10c17c/EYckwz6+FoHlQgGNRFLXyDVTyD50U28qEBnzY2d6jEDO/J/WMCe7
VIx8mp5uX/CS5xD2xUwS0S/dixHdcz8oQWxUG6x4ypsJFxwVm1v8D7cB82Qa0H3dY4ujYQP7M4cg
4+uM1qDLJtYeA5ndCVT4glYzmRv7vFq8jifAnd2lWxtjfz0S2xICvcCJJKrmSxQREy+qA1Lv6X9a
mEG2gOCVdQ0wmCSzZy1spJ57g/PcM1hknsYs6bkCXIuxYK6dkxdlq1S15j3roYlPJGenoj0YP2RT
MbsWdU2yVrwRctS7fNbWir/QjwtNshPiKmeMzVuXF6V2qTN/pvI0qjxvjTJNCMjMfOsnPS5P/cp/
XskW3podYSCnfPEH6PtIAie2aCEZV5B0sboPyJVL+HHhwCtrlEnQ5c4n0U+KpHHeX1rXNbJuItDu
aZ+a3J1uXF7+bE1K5JDMg3WPwRPZbyCwUzr+PHtYmYY2xtXKGXiSVczxH/dFXe39JQ+kMURe/+y1
hJ5ASzfX5tWdQFnoVXwF8+EY8MIKeEx1M8HRCwq7QrLSVGwCZyTRbYfqBrey2RglaZjlRCAsj/Vw
x5vi8tk/iRgfDu1XENSbuU3fXqlkvLBnMqgPrfNk48XyUhiqKBON5dFJKHfghqvFcgQvCdkOC1oe
Lf7hcAbIWG0m0oYIlV816u/F4menOrTwovUHoEyJzQmzTFIrG1A1Wzccgj0QoNbcaKnQtXeN4XwV
7U9UduPcWsgsiOV0gOIxEEc41YRlJrv9jmxqh17167pQy5EBTMyihaqwSDoq+6ghEvE24Wr9gx2T
V2JOph6UD7TT8sdsBkI0eblJCVNs5kGqnjFf9HQEEBBUk+yg5UZ7j/WJw56JsmxzldqSon+PXsG7
JeOzNihpN0QagJz1g8oVTYiPm6WNsm/Pw+fjfqxsNe4kpcLTh+QxN89PyCv/9zaVbc8b+99eXT5f
IYWwTpxebRCwh7bTUXF+EBsAtuUPrnQGSn34czDJqEdZ/nKCkVveVnEN+/DCqn0z3eAUA+9gIKIr
2YYQv8aJj8bn6H01uiMtHtS3GGf/s8bFA0h/5kJdGFbrGygN7OmQsOjZMddhcOzS1efpAW0J91zL
xYGE8JqikgCmsLfM4D34ta/uss88M0d8/IRwQR9j5ZsHMRRd98D3rn6bEwE1CsE8lkoCewPtmafa
8Zrv2hwznvr/8Ii/GQ3kGjdtikUAq5mGZ7ak5mgxev/UMpNY2OwKc7nboOewb0Qmsqo0UdsNXlwd
nwxDKXvc+asoUiuNbLVFgG+vFD2oiPpPqkspVlhYyslYOldi5M78CqlLeI9Hpg811YsCXWxGAYM4
osKNOl59zg2HYTx+wR6736sfiRtJGK0DgTPEN8BdqLMFlM1pO5prtQnSckic75f5PpB2VHW6im6l
HrF9w0PP1kIfVniOgRi+UsRRx/ACozLUZ2nxDoUvkdHc2nTMkdHR8LAymTBvYTh3UEMv4UFoM3bO
NzzuHJQyE/SOh5McDbx5zjysLyx5KF9NRa0i5TwwWmZq35wGrQ0Nk3IEgHIfgcJmF5bROPmC8RUO
XU1flaBny02LWbBoDu5Cp2MnqHMW3RXVUIvQZ6Jak7Hk12eYTBQJfZN+XHISiXKvmelLOqAfV5DT
Cs/znGFjvoXF9Tj+i/yQ5Xk9ypRslXKN9xTy01Ab4N4MOo6VMsYgQn3xjtSJ6nkiKRBhPszTS6FS
qYH3CA4qzIGUzvJ/BlwSV06VBD+YnbzaZF+yjkhQ83hh+wVHsVoxHwKOvMyiiDIBNfB9et2VcmE3
hxZH4HlIlaiAfG/hIAJtAb9sQ+2o3MuUiv79tj/lm+fizB/W8lEKwLpf/D4UEhdq438P2q+2p0NX
4ezu42occmCo2sWfYL7qaCTc8BTupw4nvyvIpd7yvvbSo3lzs+Ep3EueYAb+pHtd/K0XvUd3jv4T
5Ta8eeIzPPhMsuQGXlXoYF/tsJwhLYsQWlvz/cgW32URokIxzLriQpz6aLFaX2UPJagcPhbTC+QP
KUJ87VD2/+gtPDIGIk+ofUtvTkP+gV6kRcXUrelpWCvoXqzYTokglcXph3i9n+JyDFZmthBQXB/R
W6LeFBhjfdTw/Npqt7f5U40gaOuR6KEijBCzKe7HjZ9+vD4CN+MKOyvfsP4uuN5o6AtdtAY+pHnO
Q6Sr06FxMRET51pKFeEavej9rLcJgr0JFyxQohyPHWhE1MuLVgOMpZbrGV2GwePzhsmpH7jyC5sb
fxjYD70cbjQ6AySirKB4pat/qLJE7LKMeyUi4b2gTVGxVKIYBH8o7j1iTdO3rL5PT/DOxMcnR+P8
2FSLdMPa8xl05RRlnLT8cD8DUnUM8GkKLu/rPczWSlnheGC1p7Ymb7K8BvwTJY7V/65m5dZtt6pS
IuYfMV004FJA5Hdj2+uGpuGPn/ZtGibhQTBH88vY6AiFm3thmnXIhPa1eSe3Z1wsTWEslX+FGu4y
I+0JaBQ+AdJPzXtSWJG+xgc13bbgLp6WQG2M80pQpOaoC2NGQwo9SManCUK22yITI32Zh7r9zmxU
lteWsx8W5H6ZlGmcS6PBU58kR0xtc7ZpfLBsQw/F7/2RxgpVhF5mTvNhGwszpesLvvPqyRNlVRVI
YbCvfUWbmf5SITtJrSarehEiH2NUZ2M0IZxuQWqRJPNgIeSW4u+fnZj1lSgAM7OmkiT3w5vkAiQA
DEHaseaz2aQnKVEngNxmM95BVaiFnYW6NuaV69bWk4ReA48DdQDB29gh7kirvHxhiUWFD2KyY8jb
R2bF60KgUPZ7ZLt4CByDzIv2fzfu0YgbURpadtLOS2ekyFXcDuIaooqjkPhI2+7feh66olv2sDgv
D3H2qRTpSiIEOJJbfsTCWY3WhqpOQYU2bgdIIW2Z7oBlg1/hqJijXqMxW+GT4jk4TK83Qv6YYniW
8kUHirM7baPWg6B5l/wirkQVzMo9ZRyWthUVKXBG8HKnPazED2OI1cmLdSYDbHc/rfD18SOFX6kU
rCOKTQ1PvA6iIBs0NEmV65KARrDQCpDfHXWYy6jptqZUgQylhGOl4zkOS8el6f/+XPmHeGEwAmUB
tcCCnPaKJziTKUjbwfr/B+gpQebn8gXvHDHIo6ZUw9F1RaStlOtoFOlsOi+ruWahuTOh2whg++Bq
3eWiiYjIXK+f7rEJifSZmoCt8W8N3NtpDVTrXLrpsW8u0P0a8ix67JPZpuJhOeC7IPoblevjlr+O
kNOQlYo8RQRMn/RVY8Tsw+C34ePa7Ldc6n4Frz2Uxfs2SwCiLUXCkvHLjNBKVnRILBPaiXbcEkoK
JBGkXHOGFvIN7KxWAxtC6Tp04t+8/3yGDXUTw3W+K+eQdM81DLMU/Wf1RcikBYz/v2Uf8IQIcl2M
3Y/IR8YpWxcAvXgjA0FudNZGchYP9n+CILkfwMZcwFSnmZ5v7Jvyuh14O1c9vzrXE/HZem9U4H9k
NYZzSDQdoEIzvlfAeajn4lgmqSvSNo9fCwn7ptl+K+JQfJB9T7ko7P9FnhMYX/b/GD1XNz6eAJjl
eZGFtbz3lU7FqT9c/nT+orBdjFW9NPBkKFvPcO/BEaS4B4jlwxJoNk7bDWb7gH11eVps4yEdcZtm
LAuW5M5q8HpdI0bIzEZMY15/Rqw9h8Wta9RVExk2M2ErVH9vi6GWt13QuCyGVAofrWpWxFX2km2f
+Kr1c/uM0fj9jkD6IYFEnQohabNx2yaT/cyS3X5FpWc6WaruqnMdgRchFcxB9tpTEkD2wN2RRikD
GwTHtgzFbGYKcsT+DTSDTuE4BGhUYJQD2bueXECJjyxlkn2EXOdl9T2j4uzOWAx7BFutgdP1fAXI
MbG3kCX0/uULafRMb0E91iDKheoaYwxll75CJXNKtkaNhZSG9dgdn7VKidFFqXOLSNywbFckh0qo
4LJjscOqbdQEvuiStDBPE+Gb1YR0JxJaQhTv7wyeL4NFRLL5MWx+kD++VezKnUc+IJRE/BMBGK5y
BuJuExEn+PAn30tuC2BTwLktys+/MB5t3uCUVJMR/jmlyfSA44Lsd6EWiS13liXJUcAdDsI6g9xX
JBL2KUbRJ8co7MiLNRF47u+mpSC38cvsZRwdEH5LlEnPia5bj9/tmpOKYwQPzHTji4dVt7t1VJwz
RuweKPNWfSleJLFHIVO3qj3QbZgW1+j/dc5bE5Ya0z4KxfJWqw2l0EHfbi5XCk0fO4MRXFLg+Hth
BLnt2gwS92tapf9yHSRFcRbAJU2l0po0OQBYq2ltNq9g/TNlGE51ILubpRk1O7PEZNfNYfboPGTs
03nG5JbNgLtTNPNuDnbQUfxdXgFO0RqkF2mwk46grkvP1X4mb6wskfyUUQhHYOR23OnUqkNsrukY
Amdl7eYCEAUr+EOPGNVGZmxU5SEA7NUvcnlG56FvwZjmCtIw8ddMYudsHqoU0IJe7jkqPLmX7qs+
XlEVrEFJX66U9eBauR7sIdH3PyxTjsLc7+ykeWW6crD3n4bnCOVBlwGXqou3vWT9U7RIGG7CkAR7
mmy6vUKW7jJYhavcfXWcWoGcZGm5+i0TVM+Pbakc0zgApB1WDEWAtDZvagjWPi0zfh3yOlxd+Crz
PKaZ16k8/ieLOda2mf0/4LYfyUNqOjG0JyvUW51+t9IUY8YD269tSirZoZAnJ84/iGitNRYHX3AM
vnf6Oqo1APXLxMAQLFf+Vf2u06d3RLhp0VrkDuM3Y9uZUz/gWoOFzndVgNoVz/a7i0aLqGF0VElY
ipq7/bToBhBzR3c1MzVT+z+3io58m/5HGDxV/99DJfeVYul1cjQiwyxTCNMVKLvKNJ0mz8oU2bQQ
qPcIH3HsOhmNylgdWssirt4pGbpCIQ3n7AsN205rviMDselHVbEeXOFPsKqAWyCcTpQTsl3orPcb
PvSrJZz4PP844Q8fvQ04DnXDsItTf86m+5qyH68JHKuBFQjdgPrCN3C/qRB88jtcA046mmx6/58r
tPr2WGJrNSQwN1gKHSOHhK1M/TafocUXwfXmcshmO/NsrWW34QHQ9cLq3i7/CpsNBzy5Rkp3SATf
OJFwEtfuiihL9kLBA2AmV+6LsS0S7KW7rRP4YXvZABbhTObmUR9kIBUL5nIrCBrg+cUbkCNCwuEv
M4pQlAlul1qovzslW7GL8sHzAsAkFVfMLcKty9gAwlJGPsC5VheAPOLhuQPqz80cB4McM2q1L5PR
WxXCM4SA4QDSDUW0msUq6hKPYTp5lT+kPupKRVcMiGNXunU6+LiPL9cj+KevMSpYVPCt0XMhKz+w
cKFM9Fh+dXhaByEhLly59lqDo52rTa3ZY18XHDiMRnAn1zRhEKgduLbIPoPezj11V6PitQmeb4nh
6WF2P83jOu8jrE4CfO6q11qQqeQ5nchdgOzQl8OUjYaPi66KkWu7e4IXMmVdEAfoLKdM5TkRm07u
YlK67SlkPFxa2C+OrqQATBuXcboIVj2SKLCjvEevquJd27KtmKZwAoCX3XuVze4LTluzrgiXblct
1QSbUQStuF4maEXqaFvk5roZGAbqWAjF6bsp3xeKq75dxRLMUvKRtRssLYZ76z0Or3Nt/nwvGo+i
yzYwZHM2iKA8nc7dx9JHTutNPhBgALSeLZ6GovU9cH6hz6vlTEJ5S8vAi5jt7d8cnczZJrOSzlIs
uf16Wo6kCUB11y2Fh1g/5qmL17+owWkhxAYkYrhH4qyS+UR5I8QGkVQwuQAfGk8vglVKiAldIAuv
Cimi6d8hsVks8Zpv3N9R/xrcRYck7KpxcfMgGodNfmXt1qhOqKJxoKtAQj9r2pXI0NwOGIR3Lkpa
QnJYCEYvIzuOOXSlHBMenr++ZDFLY72izFYLK9F8y1w+hp2MHhHdMiBu52xV40IGBfgcPdTEbz9q
TPaXKMtVjecUaqMNeCO6nx4Yeld40YAoNSYzWAK0ZYLPS8JxIC1Vn5shEOhuZmpRGi523MKrIpiF
foy43ugAKsZxVZimR08Bp/b07gshuvzBo+66+h9IU4fKuNE+zCXNEAhBOpYoDbvU46XQ7Nn0IrCa
NHXmVr2fttmLW5h2x+0UogjTWYNNmiyWBamV1uVqHWcJcsmAf7djcVCIpFNsvrdyq81CkDFndJQK
o4Tk1Qq3Uw6hGLam8+rMrF1V4ypvoU3A/JimN744pZ3ONINs93/8Mcv5Nr7LJNNy88h6HhhQeNTb
h0pIN+O+LicFl2hhgY91sl//UCj4fzC7wAX87YLPveq5zak8VnodzXusYSRe0ozORhAt8Bip0bSO
mm/T4vfNwgYd5uAsrpXXqP/OqjMFY8SdzyjdNhAivY5nI2tS7222E/E+BCjbcQDdGiM++Uvgkjlf
au6XDPYPT8gLY0cMWA2rSwMhPv+xY4uLmjtKqryKweFwsHravZ4QFST9/HqyEmyr1yaUbRQOjZhh
heUuRv2n6maSNZfvK9kSTPLxX2phyOSrwwPLKkFG4X2MGJw206AtEr2ZIcbh5LcqXVDFY7rCSptQ
PcHp7/kBOALTnhH6KmToNyM4jPu+JMrCYJt6qH6YoLQegBab2X281r2321qLho8MWBs7DwhPIfjQ
alpnt83cmbg0OhcbKsYMWc3O5ZF4zdC1e4c1MRDByk1OTlZkv86HYhfBRAL8IJGfD52zZs5XavLp
KPW32X8t0vQkQDgO3cCrQTI1pJ1kdgIBOBFsDAvHdYkXLRLKkdl7k93mTzDYFVTfPlfj2O2bzZnh
0WjFZciAIXfgeDOVvc74gAPXzAG1e7tNSDXsVhq7FmZRN3Cr7TjB+l9xlHrq0wy0W/3BG99MA7pW
z2bZMRLxKp4HfrQzkfkAf+0gvfAl4b1VX/WDLpZkgehjB9qUgeNuR1cbpRtZEX6278e7Yinw5BKw
4NdqVSjOWf3u/vNqYUjngT+FZJ64nyUzj0tBhykgda2LztP9Wh7+wChb3KrxpREkw6pZhPMpC0pf
NFo089Py6yBE9V0RSMeCQv6RzzwW5zvnCuVPjN9eVszQ3yHphA13M4zC3LbPbXGDUuAvrzBx7vQW
hVj82NCsVFsqOXxrhOuDaDEX36KoB4ncEyo5/HFmjuk6yTJ9Fsq3XRkn+cf/ULlh0WAuqDXI4civ
H7Nw+CCKTKH+KHYaEnn5l9bb/c4aPfV8VKnOLumogTU/4aKJk2lgEqdBvotvozGNI4sYUgS6ga9n
gpw2KssHYFij0szkFzFKvMzQqHfqL91cooL4v0HYhV7GC6gJREybHged7BwJLu68eHXq594rgHTU
TH1eJngbksVypvXBR+Bdf6XOu/JUt1Ym2JPBSayDShRzeg8cUQkApvzyh5OYcU5lPwh//IfN9QfZ
piN0nQqTO7PJPgGltdj+5VkPuQhE7nRywNyqQzoahM8sRxY99341uVmW6ld/KqCIc8xq93xOpO26
s73Rd1BIOAOC7NL8cK1POZ+dRMwAOiqezGYHBY6JO+pstmJYoiLXFPNPZ1rX6ANTS9y0EFzhWuHT
AWm/c7OR+je4BhwRk9WB2bAtxi9FnSfimyfzSkJmkTcRdvvXfgfHP2dKy0JcbDDlyWbut66aD7O2
/X+yUW3O8JChjbirZzWuVb27xznq9bJZZKqODPxBllbYgghm0/phYXpPfgxL1XnuTdrvht95O4/d
Wh5zmcb7e8ePuVxIwfPO1u+p/8PrK+r8p9yWgwMAZr7P1k3wOCAGuLR4xJT/1S7uYKwdXI/WWqMy
mVCB9EK19E9/KgtTtmmLtPqtecL1iFDgZC3X7JEiG9ZxdlMVrSkrD2bnnPuIuIozSwE7E+v9V65m
rXcHXzBoaZgDnIaYkbrb8vJTtp9pEqCLPDo1XoHTN7WeNXsMqN4myjpbmJwC4TbwuZifIi8q00Kl
+bGWssAVn0nTjPM+EbfdeaJwfz1tvgzFnkbWYQ/9bw5TzlifAE0tF49DAWn90ZkqiSGn/rHYSqRL
E5hDRT0XiiZVQeZhUL8AZfO77IfIvMxufhvTqHHDNJAzaAXksdyi43s1CG8KcFh9hsWOcT/5yuzP
vA6AMd0Vwda2vDUx3y/CFMk6bTKmIb/a9+VVbeNk/CtSLpFltRufPiTaOr0qHMnoQ088cIQzBkx8
hsK5BQ+YB0sIHbY/siEj49/SV9XnpmXWgm6wNt43Hjcd3+CT+hjbIwNspF8EnCDQyl/IL1O7EGma
+8U981nec99KcLwb78uPud6SQ1G7SOrWi5mWD8v1A+Ckp0gTFUIceF9X2RCQ66zISKj8s/PN0kC6
U110djeUmJdAujL9okmafmh7MIWpilBWmDW4OCBncMbTFk4esPBiFB/+EKz/3ZMWubxe9ufMx41o
wFq8pWFgC5VYT4Ciy8YvVV4GuewEUACzQiJU3MC61QLrWh/aO8lkRAk0zw1AtBmQfzWJmRJqWca9
ME3J+7wMOdgOzq9NDoU5V74qShtwT5T/S6qjqbAruKR+QyGzNKfRKiHPPtGOYVu43FFsdTJGuAEJ
xEPGMTQvc6pArmN/BiPUDXS6gbvI8A3gvJgaXeHdNoipiZNuWvfhfgSPt45eG1L25focT7cAG65n
EAny2LFFMvaTSaTmoj1psUoVG1gWdy39mW+KZ60xdxZBa0Eu1UuUf/tDcIiIjvfl5jMBG6xzwJ+g
fiFC1JDUebyPURjA9mMTHOsWotddIzPvTv6E3b+tYVI6zmDp2+ChLmmAC7rbG5tUeRiir7D47lHj
8vcjo54G6URx455+WkUXvcBWJeDxR+nmQKo3XWxny8TG7r8CfJSuoMdraiCTt6n4qhTMBkX7SHpx
T0imFNOQPYQ01nHmMYuZvykuAqDBDaqbrNCH+stwlxxFUt3Kk29b2uCF9aS5O0HNQNWEjL+ii9wI
p0pY1LIZVY4JC8ZU1l6QO+G/+ZQKALWD4G51B02bgtxFO0zP9F2uu8k59DRY/jwxjUGsL4/F8A0U
z/mPIvXUshKqfrFr4BbFKvBoRQdjDHgvkEe43t2+fVlNLhhKgybxAIdmxA9B5839Nr5l4mGoV+na
XBIciFw08niGnkg2qerSJXX3QRKqNiw95Aa5Rj5Y8eXRMyBpoDgkADbCFWxRxUIwTpUk0ibLQfoh
ea15e+rCMzX4vnSoJG9AH+DxWGUW2vS7BRI3t54Vhku4MnH0P3MFoE3kHxs7/02PoYKvyv6gMzRK
vRI7K7XRe9ING5uKDAmqbcCzS8AsjRQ65fHxttGowmHb9Bou1yrIlN9kngKMF894piEUAKYz6QIC
+UdKIE8mCY3kJk1KETrhjFYuCiJD/ZUAEgNaPw0K1g0rTGtuwy/E6Gamu+cr0rFeEvYVEKC18x2E
WEjXreMcPaz7ooYKUN1Xbi4hXmmG2qUNxIoXoAhIga7UuRgUlVs4XNw9isYMp47PQsuQojYBgzLm
cr+CZm+B7OHnSZyhsVcmE9EkO8bEzZ1Fs0ta+Wr/ZDT0SVb5AtaiReoknYQ/hQimTnY/YYxXVeTh
cc+FvIvbZW02ogICjTd+BtPFW4ewz9xliprv13c34jev8U1HlWCnWpCQCIn+UFeOeQY2rtztNaaB
EuhlccwBu2KEil6e8+YBD3u95rT+7crDyPK9ScfumsWs45A5yHH9NvFiVJEpdX2zzebTRiZlpZA8
JXMwM9QAty3LtLMmdoOqGBx9OEs/UhSSnYv8QwrcIE+V87bzRy1L9RCLqCucK9Wcfku+yG7Qa8B+
OOBwOKtG5LRPHOeugJOiwkq3t/JaX8jTpT205WqUVTrOxo6rtguAQqqNipmMUEMJAH1vlYpBXjjd
1k8VBQRD854A5DFz9Lo9JwzlVMy+Bd6Xs8rrvS0ln7lyvjNWKWCEju3piBJDVgkYlN3+w3jMpJCo
shcnmdlRfYJ+zu6DjiRf3QRS+xP7d+7OhT6CatWVAqPxwTt3YoohLgYJj9b3dv77z+Ohas4kYNme
kZWCV+1mg39sNtSWBmmXJp5d0mhaDlvQS4fGR0KkQmRrmyOdo7aYZNt+z8+Wj+5Ms36tPOTT+zfW
CCugcUWBYtbTg2K4L2UE3GHpm57cCsrATEiKF1/07F4yNX8SrEyDoJP+0xi/J3kF1q3H9v8fZArR
s3LkNKLYE4sTbfQDvJ6wTmfi3QogNO8xvHqFjbQowSo/2tSUSNXW/tCOLI1vPQBB080KM+9cpmJb
K9VPA54pMfUo/JTZm2MVR/QFmyOw7uvz1kS0GHDGvC254YasbkIJlNzbKoET5hgTN74PQ75UV8K3
yAAFjEhmgcHRolXOodvkvqVzPU2Arvdw2ARMfXLDgtiLeMZXFnfa8l0sMSnJGMrqMn4KFNvg4dmg
tVRPA41SX/tvsWEyjb6WagOKH53Q3yuSyiI80L7baZ3PDlQU0ioHyF2spkO1kD38nlxXwCFNV3xf
2NPTg9kyHuZIo7Nsz2e4Eqjjl1kL5Ie/tZTn9ijhguZHRy0HzysaUchQLRzviBXkQZDcFin3so0N
XgA3SX6MzlOYALwYMYvurhuuv5cYNOqFwmNP8sRojYiNXykXOUhurUMFsH+6hgYtR9LVLnLcQzjx
AK1SLnRZCzSEdubjNDjGLLraV8gQSm28Mu5V4Sks9CPp2kfB71uh8A+HHs1CKHIQKm4f0w28tNuK
ONzuQ8E6335Cu5/HNsfinuczxhTaqey2Ew0iExXsT+ILvRLrDnryPKUjwZfl7VyauQJZE1VkpaXO
TuQX30gOcFKa4feFo7cXz61l4hQy93j3ezpK+csQo19+fHEvk1N3qGDvG4iiV3PGTSoXPBuobZsO
iGeWm/OjS23+b4nZetBAXfU6QZZIETkC7KtDLTj1U2MOhOV+QXvM3TzU7fj3sHTK96DIdCVjLwLD
MNz3to8Jo5paiA+Qq8Rr84dI8W3cU0vo1FHvCTvGOd7UWlNNL88n1p2upMHGhJqqbnRFmOr09mT8
1kFIp3r5YaJEZYNtTcJWVhVT+KUXOAL6VDipNHE1MXWwcweYyyxygtT29Nv0AAmf9OjgIuMR3HuG
5V17xBl+RpiS9VeZV0wKfZJuOK6t6jh8eYO+9QJ07CkGlNLqaup6q8gJMAu8jVZu0m2fI7dv0LlR
FX0A4ZlUCukbIigZ2p32I7eFDnMyyWGmj32JNJDEbV/nm14mZpbXCY5Wn40seDTRlqT1KzBIFhGU
J73cY9zbtnKOoOtHKlkomh6JtpaILiAZUp9OovqRzc1MmVJ57dOzEERhGyq6+KclID0qPH3W9mbA
7lagGm8u8NCLnFLXJy9mjXhDvdFOmjz3Lox8q1F5l/u45CuDzN7rCaHzSw05Y2HSuC8B9z6ZOnO4
NP6abBSpPEG4fIz70I2EQmLHIlECgSeDcL5guxB06fBjZjNYJpxGi6VfdeW6I7et5f2A7sF6u5cC
xBIhfpO8vXP+Fw2tCT4vV0//5VCUbXJI1qGGeb1CrztykjnILrhDY7H+3jOL6cAzxK9EoTbTYM4g
GwjANignbThr1i/3liUsD8xDUSmRFlqbVucdYfVhtiqLwHt2/yr7dtIVvVFCj1smKdhX1cdauq7/
zBQOriAeRqJMGo/Ag0gKABBgSdj3akYZ9GbtdDoId/Rj3ypC/GXwCwaRPjOrL8PaOBjxG4uixaYD
FCXSQ5j+9gmNbheICbhAUFeXVVxrSZU+cq4TtcN1o1XjJRjElfy3MvOHtg0XdWpECZUwfS1RgCuM
fqQAIWbDERdVkxvnW/Vxbp92p4r5lZ4h97vAC/s3qNK7abMg/M4f/TvhnGydeBOH1yfBGGpi3/x2
mq5iqw103nHdg7FhTraaTaKET8gO88PteSyiTxQNC73ptAlxMVx0i8QrxaF0/pblzoiDxnpTDMlT
zJRZvUFdEcVaAjD4s2Yuarkyr+ZebOvJUKrIpHMDc/Z6yIAfuO/1RD0IKNF+Zq6fyfJ/C7r8ESWO
VpcXZB1v9/iC8drzX20atds9B2sBt80cIeuuc9+LGxyUptbSwDbYjFONVD7lsZi8KOKt3Kemimep
uZGP54oJv6pxNEvOzXv2+ofTBqcVZZRdOZxVV6NfQZBofhqGlqmxkHT2E+UpNGn8Qix31oyz0WFx
W9V9CRbiOwOeiOYidrFtLhciZQGFGSTkXSPz3BYId90+j2fXEryBrbB7YzyXfKVCyJp+KOOzcGb0
d0jGQB4ozZS3inDOB0HdqKiNOCoNu5N617dXsiYK1rmH8XExHUW8lmJdRDiFVGN/n2OCOtUin3pk
mFffoKFzwxJtv9KIYioMBdnmDsDBdJy9UUqTtp1hMoBGqNA9WQrTduCkYdNs1QFL1H/cDI2yHPks
lqR6oZomngTRlbuCNb5piNE8bSFVbblLUT7Z+Qmwes0s/bGEJYsOUVOnXlVjieSRGA/+YoiSZtAd
BxzN+vDyHQcI14TEqDf5reqruzOMshAU7owcgU9k/cFiGz5Sx+GQnfCXOIHmzjeh7IfSe5+3eK5/
1Qm7qYQLxDunaEYW/7786NEf5/dN9gs9UC0EQZQaPMqGagVKpLlOfmyqB25uziAponyJowksmArN
eU6UYyFxSPFU/uWGiml6WCB3cbcwKvAavfKbWR0VHfqV83wi3W9ajoUL4hlA6mhNkizwXFNj6W41
1ceIKiFtdLZOGNcV3+SD9vcldn64Up2c9U41kRiSgxXka8qmsuXm5Aimcg7HlDfylFnvaNUs39f9
No+lADhaQKPEh95k0JvkkG+K5PRTs2ffqMIrxOE8NOpiJ3Ygwo4gsV2tRVEOoWw0MRb+YRRTivL/
uso0KK2epaP8RRpS04L/68zvRt1m+r9LZIvqogSTi1BSZCN45eVjw07YXghMeKPasWx73sGZMJOW
LcHAQ6uEOK70xIRsz4/Bh12XNo0wlyCOExFVibnKJyFCaCzAcxTvafti3RIZpcY5lyMsOKifgEA3
xZRKD143w6P64azEtKY0xwFJxEdwZUCkfyavZpHAQhVFFvQ+xv403c4NQsi3qRSzUZRrhBUU4ZRX
j7P57wqeP1vtgChsQ41Q5p97fNIo0UQCy5zSNw39WF7EzF3VVbiFFvIsSKinZmCLWSOncztOnOEP
4HaAtDiMgSJ059iOwcitRmyFwmLQZpRXjjOvDyHh5m/B7MvywG18LoaJT9mGDEmVDprq0QeeTNbj
Us6sYKHkBsiCNoYbmFw8H1s7nw8x3kz2dDvqAEpQrO0kg8jQfU6ShWljXbJaBKymgzJKCIaXUTCh
8jNu5jxkBfvjRi4gJJGuz/OvNBlhHmuoSQq9ZqP9neEcgSKwX58YE1ih5Vi4aq4p4NKE9dgJO5mS
ousygSlnexIJmvOvqoTXtvr1qskOikh5iHeqkxbg5FenFKM+E/iZpFmdRX5u+yDpN/56MPU7VBpC
GN1L3xPpvMm+0Zr+SIRoG4EVqGlCL9v3XwmBCAqxaFFALDFuSvT6tmjU7Pg13YYg8UkYLMxWGQuE
+JH0CbSAa6G9B0sP2tSmDVd0mXL+M/XnMNFk0KtQx9GrLs05OrSPizp1DVkOeWDoFPMcVe5oiV5z
GHJ6ZC+C+gLui1pZusYHmezCMnDEkkj/2hdn72kWHNTw6ceIHqBn+utSgHMT7OBUGeHAE7J/5OjH
ryVzkBpTq+jKCknJUFj22JXOu4xUYfMvXWLSDq6dIr5piQoyNZkhn/rJsU9OqBzKsTx7vBfrq1y6
j6LBkHpwXkAoRaWlU+J06IBZ9SDkLf8hLlJDKDuYm74RyTfxR4hRsxMxQPC0mFtf5jMJ55vR4Kt2
LwrZjRYtPGyBWNfhJu6BLjV2HIOuIbt/Gb5tmwDGIgMdmMJO7sec/723j/8HeaMuBKUiYqscocTz
igCcK0dTJqWXfErM2dz3nK6zsnoshfzpvsVvjtjYLYRDBnJSj1WAkWMfS8Ur25zEG7exnYUfnfyS
XANQknA7xI2EVp/KfTI4USmqA59ZxYk9fsKFaxOf0mds3DXj1/KCAY06dEP8n9wWXHgZHR700vTU
lpQ/OHKYuHIw7jLxbz9ZChjW0+CerB410RFiw6ZLbUgel08BWIK9A23Trp9i3e40WwxRyFnvwwo5
r26qe6Oyr3wKJFnjxpOBQfeHPr4RgdKmdsIj/tbPExs5diuFbBf6kekTM8NpfnZF9UWqbRw6+YzY
UNEEZVoVD8YuPvXtvARbVIzgYMkYm/b5zSv1c0hHEGjcEZlaa27pTgkQSWAq3/mAiyNJUtY6jdZA
Us4HR+v2wbgCT1S4Q4IJjb5LC5Ub8w/iMgwRurnyIG9imO7xnsNt7T+mFLTr08FJePG78QKoeaTW
6mtHwkxhacQ7f4XOvWyq/LCMR1baz2QDUG8v9nl5VFhh7xPOx66X7DCGPw2Z+yzYQgmriGxBCbQ7
ruW7FQGrN4oOFFxp7njnPtJsa2BOIY0CPxe59tq78UJ8qB1JUGv91x/QzWKrxNnHmYP5sdDYtR3g
+v7789GmiYJQ65zWScB2OHSce9NmShtlRKdKzVUJCtKfVk3hgDzGzLnduWir2jW2E5ku42MOqgLc
TFi5YDyZkLHctO1zCus4WlOdq1qsvfIKU34yoDgt+GS3IovtUprM049o0LDAHXizTA0xKV8O+92/
swXKPtLOJxonjVkf4IjxMIM+ugo4NIGfTx+bE+StXcVxlioIGjV/EegJM3VbrT2HvlXukzH/CAnS
fP/BFmkXSxgG29+zvnlkrFbLpqRYWrR5TvyCTmNTqLRtl7PwgLJ2iNDuC04hTrL+ZqSI2LKUaTSS
wYLhcRTos4qH5R0NHzluouSuMafpu5tvQqW1BP7bwN6Wibsswz5dhV9gvpOtD1Zp0I9TOXhdGnGW
QeCmGgLmuokYzUr3jZGUWMA2fv3lTBaMmxFVlTwQSUuduV44cVurisugJ6E/TkwNDbHAqGXLpPRZ
W+FTZo9jQ9M6JPRqYUB3e6M1djz+saaVvycOY5z+LMV3PO1KWAzIrKxVRn7z1OZ+nXBZ17mb0ZCK
EEJpNAUile4wmqIe09iOHN9ss0z4cKwczbPhUA/lB807cPqDJotEdAJQFBXKTcwkmGIk3tTuRjNG
e0iPPJorJc77WmUba3MO/8zrkFXaarCKBSUtnQbM+PEd1csi5zec3QZ4JAY4kLlnDrWPVwL++yY7
ahqd9K5ZB1O/U8d3qb3/0BEk13ttExnJaRVw+YQJWRxcs7S3pBazKKZbRDFR8cb3CSU+4w4/Ckwh
Ub4yYqvGMXH/GBhjhUeo2gKQqymE36GflmgHyPbP1SDIRGKhyY+CGdB50qu87BrHbM9yKjMwH1Ky
APKPI63t6X7rlM6UpSEpgPiQCDX0Ite7zIJ7gm0OUVlSme55jcDqOcq0Lq+N3kQZ1KCE4/3Zsfjk
WT83e21yXnsDVtNLSJR5CtDdvW7us56wDHw82uzR4e4EvLIDJCGei8aRKqPiR7C78WDRcguoyX4Y
7stB2fztcDVrqDiXZWFfiAKiMDmGJyAPeE2CN6J+2pncuBimdQo0tPRIU/Iv2wtUVNfYphNgRXRY
hp+Eh82qSTfeg54G0PEoQHXU2PF9lDyrSps9xt6q0s/js2zKOc9l9c5+yOH1aOAxWHX+Iw62+uN/
tQ+o5HutCm+TswFL1f1YNbF3ggLojp772dPeGJesAQLN5fyNuvlw0vjY32oQHuc5Ql2O49idK4bX
js1Jea+2sofI9pPFxOwZneOVPHiAg9nfC4An7DCnvYCWleoGO57GwMU3Uf4z+y+kZVFOzLdI3FbB
AZ2uY/Lrkgb0kVGPFCnpO5ni1d3A9Dy8/WXo9KlSLr0FmIJ0azoMsJ2OgCuuMy1iNa49P4AAefYC
WWwFlwAv7Qj/Pdo6t7vU5hoEN2T68AFM7hlp7ksLzUbEeoSCygatTH6lp3AIFDIjHcs8se9yNNKN
oD6a/Ew4Ym01vgdEDkQvA+rCTOSokKryHuBtDYNgiG4jWYjRSpbAcbqdN8FM919Kalh7RUFhJFIL
8GmJfKYZ+q4JtvpmJW7jJa9NU2ByA7ajxjyCtow9+lMoeGbj3I1GaMZtFb1O5WN7V88tiWCP5QsU
y3hd8g2Wlw1VnLib3FHl/mAirIMWHN9E7cShvgTC7QxXRP1rRh8of2OFcIkjOYhAUPyoCcXO49iK
MYafkPjZFZOYhA2G5pAPl6fjZvAuCgJpQcHWwhycBXDvDp3//2jCV+c7qqI83AcDoGoMsSXAM2db
7aMYgEJLVYsMiYY/RteOF0hrjAXuVuPDpJD6fnjk0N3g6m168rIEyVhIQvllaN42RG3sssGOBSIt
pgMafSQ90n9RNqT1ZG2Z13ZWEY0HCSOdH+GWmrAkCM2QysH6iHhNmdA+9CNL33/w5mjd4NeOit9M
WXlZBI8RYovtP68FLR07nn22fItkTszCkTH+Y4lBihS00NTjtE9G0pPZWoKQ+ggCb0+hZzq0xOtm
U9uLP85Mmd+7UeOfeXI7slb4LPo1gKbjL/OQOrOcY/jktX4w8G499VBaq2O71QzSK46bP47W2FAd
dhl2mde+3TeJggnw4yF/bgc9DVY7M5sEgxDTqsMxSOyLIN3VP5X+lYTBrY9XUc+0dNqIl1aigVpN
L28dk0dHKCyyp67mWW5wfYm2ZqAFTFBSx7sUiiXLzV6+3vrQsOMM/ScuhPGtQR9X9IwYxfcMpnoY
EV1PYzDLUgUdMufoQA4YNeHYM6qB86C1YKoXZMGDou9OCUeJ21pRKQ71i6Lqf5U33/5naiPHBvKg
oIU99MKUyKcUUQqNo0H1mGOwkjXFKU0E6DXVZFjiNJMFr84yOxRTLfLWe2ASpwZYp5orlO060PBW
MquI3wYbxZrUrTYJET9xpEXIwAjB7+hDHsCT3Dts82aDNYxtz02hqUZZBTQGSOTDoRdEZI7euhQ8
zujEwAsnUQ/OUT1ZLhc1ielY/FwdCD+BtwUnRV8261V4sgg3Q+Cr3lp3lQsJgnXJtQTmI8vLSTnj
ocBhL8fb0RFBI7LWdVl8eTYYz+fE7efDN6r4IyNyHGPIlxhi6y5OD+XOsOVZKXSKTMNhpYcsGdt4
eIP5TRwv0VIF9y5mKh6M7T+4xsLgiCqgNfP40cD2M+aOPVfvBC/tyG+daX54BbVCBRKXX/MzNUuC
d/9dehHYEiynrVbAGt+XrKd+ebtbwjMamNGf9IZExYSr9lGWrEFA4v++q0CFRsVOFC78Mw1+JMLg
wdtGSX05QVEMIHeMdqSkzbVSs2CCBaOoxgpjIpjKIy804MMBQaRw+i127KdTvqkZL6uzqko61UtE
0vc+PDvTD0lW++detiEmEnmfTYPLD2xyGHmrkA/R9N32Zw5bpTFQMCXcLvsf5fZ2TmlWChGhPcPB
P3GMSDzAFO9TPCZjxcAzco/w0lUBreylmOrPcwuml9Pay5tsAMp9shemd/J3owWPRr+Y0bQdfKJX
pssYoZoJBAqm1l+YLiN/R5gBrzWjieeTxpwuHGF4oIzcAuovSqJNPOnzbr3ia4eJDO+DD8XfT79C
JYC5jjQePCD2muWK8xFocNBTG8Rwnqzeqxevblq2/MVfSCqoGw5wSVfYWCNKnJ8OZpNodY4Drs0y
kpmySlKI9Ptp1Ev3ZbyHkcLvn5s3scaanPB5DWH/XtUuI3zejFA8WXj4VThr36qm6/UCLpsQu/qa
pykojN7Y2hykA3CzzV+9BZhgA5r7cXvSyEei9Q0IHyJ6nJJA2mSTRJbolQ2oLMlyCZmKgWGYpRmx
P+7JNtBrvKPkzSh4+Az/yjvjgkxyAuyoNx1/HppvYy/YmPbPnbPD3kC3n7CNREk/+9X6eLNQ2nrF
a3c6IaqGIs3hrS4IHaAAKpet16/hMCHEa1oVCmK3f4rkkSmFRjhjMqPGtlST3Oscz61CakUAp7gc
LkB5koNeK66jyZWNemKA95PenrAAaA+dbUzQGqOBhUeo3nanDsajVoAHFv9lmQsA3Xo+CTeMGwVt
TjRvEwE6cdZj8Pmp8aoCTCTnnGWSKstXN4KSeoH4CchFu5wrWGIo6CCZKzj+zTrRr51dFMZPg5zv
TddXt/Tf6xf6xnbj6esFU9EjOBzy7BDNmSF0bL2skabM4kWvpnfTjKsYPDDJoJSC2V1Qf0LW2djl
emTz4QTHtxV90c5TJCBJwndYFFrQg3hMoTFmpq7tlZ3PV8NBoCrNNdlqIJeW0ISliAizcqUcP8kl
9+KSbOu+8bmwvFcNQm0Lw9iBaR8CObahfYIaF/9BN4LWgeAkghaLIz7BRjuyuyULlHj9rYga2Ipu
Ot5Jcxd+KAUFE2IE4IPRrRFCxps4a5d32aK/q/VJGjRIsCCefN97jRiy4jMuoPY6hXfYQ+QRFaLz
CqSwjcBQbpF7eILqfsPLPAhVGXt0d6F5ylaNivuAmwLXzKRXmGfIiDjPuAjGa9eOGexD+dxZIfIZ
JBcc/yZgy/mXsAAFuFg3Vbc6E+QWiyj5bNptJJ6PJsP03P5LgD7cKb76X6oIC200RshV/0U11T90
oc4E+DSEHUtjKoOPMdYvt4MQAaRzpsvNVeqyJI/h8X+KSy13pDQ/2zeN+PjCUqekbaS/tZslOwSc
kvTpn+1JxUd3MJEvsJpExTidC7GjvUX4+E5EP20EVZNQFCdxCcThqcpBz7bEYnjmEN0x08QWwY3X
hTfE1E1aqHQTvBsZVmPWnaVR5qwHFct5JRZyWCOeg4DNz/Y/gPeIEBSl+vn7SU+DE7sepY9/rkM9
a1YZpG+W4ucV+2aC5WN1Y1vsuBQ+Eb6KcHZdlxcvkYwnsfXHJ1IVBm5/v7/ha81FdKgP7SGQTdJz
PT+0ndZ5mlRF27Q4mp3wny/OGL4OYTb7IRPFwoahI+HzQU+2WeILdGWWobdA6kBJl3Y8ObmLqLiJ
4HJiL5ZlqPvMXPcwife9OlYM8F+p/1OGmu5Vp8h8GZ41xGX5Xv5y0l6U6UouwoPDsPWq3YyupY1n
VxU0oUOWZ+j1a8NQDyZfPkc8LDFU6G2edqFxBBU4HT7l6u2G3TZO6iGuJakSCusPMk1E+h5VI2q0
TN656jU4UbsAAlKd668Bu+zJCqysqAb+AOv1ANMCatIaC6LatZtOSYQPzJHVnFkaarLRHMAxkd1j
0JTTP4JkOT4rbr1GJgSIQVyC7eqzQHIwKQkbg1naOaGh4aoUYXAm+w5uPuxgSNgR45mzPAsDER+I
Q+f+j4igvFv1+BEi9HOqAnM7OT90kmZQpYDgStrEcvmoOMCejsOYjSXlJRSLwnBvOCcNSOH9K18T
w2BFH5xon/CT3VpvLAhej3mHw+8puoZRIgQQ//W0CjtMe4gKWmqDkdzRR0btrNykLYz0RNQh6Quk
crA/y4C6HgnQPqtWPhgnsGO8g/YotvUayngAbznhewVNp08N9/s8S/ofPbR7y/lGnnP666rjOXsL
ksyXBr92Dl5boyWi6scU3ccm3/wScrZLBiQJ2jTQp3mlOO4b6DJ8CGN06GYvTZl2oq8YIU1MBm1l
T3sQdbnEtP+XqVqa2zDAqR5VFx6jRxmMKL0n/NS7rvw5r5TGbR8Y/H6WTjy1LaP4Hv7xzZNasC8O
BYXdsOV7eoRxteUtb3p1WKJpJJv/7hNNYCyEbewc7f5sCsQPSL+J4Od+S4yqG+ZR35Hu9yGN0ftf
I5T/Z/GFSR/ZkaDHBKiI8HbcHsgntr1iL8GMWd/1veZcmUtT4S5gkDD9Zqq0ibw9m5VPy/N/io4W
tYux9l6ffLKkTv1FL23PBbgDwQQE4Whj+1c1eUg0UcoXixnrfqFCcumkbPVaZlMQHsBw4RkF+vG8
85jJMG5r8pK3Vbmj4MtzeKs4cGpIljHKaZZVwcBFMfW70CdyBCmXwYMO75UL8zdNgea7bpzkvQeU
A8IywonO5d0pBi0kY2PdCE45YG9PfdYP+7MUREa6N/KlDg83Y0is4TrWV2Pfq4Y6jYiItjOkoUZP
dLEcg9vUsbJduMsbiMNwV5Swhh21C3Kkh1bI8P9tRgTXKUgxjW/LyqRCt9XAcM7TgQUZDZwABWoB
vC+k93mwx+LQ3Upf2AjOMl4eYhxl0Cg47oalBBvCSouUbBvGO+tCdQEKUhbW9hY2ZaZ2ydXMLjrf
UjcWKJq1/ACuTEmSqK0uh7vXTwhozViKlEmBm9hkfwctQG3e2nTyJA4rddBOT/J17kFl9F0+hiYy
Ek9+A2DoP5HwM+Mj6D78RyaGs5XDgTu30jnYxXn8j+3hF4PnHpLXxFkto+ZdVkziOHslTa9y8ios
gYKCOEngaFuU7mdBIx2W+N/jGeMPwczsHvSsPVIGhCNe29QpAxj2O6ZjuA5PG5JaAwzj0YAFIx+L
HUSYfvvSfFgVsXeFLoAqbBwdyQf8ZLjjuxq8DoyqoPAuTlqlS49lifDmjf8LNAyeQXd13ocyzQUv
w/PjLnQMTQJriJx1QmDiQkaXov4pSv60nX9dBex7js+ksm7DSuvO+KfncRW4kEoaakfVcntRaF3S
W1PNywZKrmLLWlYqoLYyfsy7VToyG10kB4fVGTIBQAKfiiifprLuiPyBvig1++2BCVM5Xso9Nmmx
s1C1aPn7NNEnVg5Sxk/UCTJMBXGDSX4pJOMptz/cxgrn5I4Itt6KcM46/JIJL3+WCQvB8uUYHwdw
/gfOh5Eyjt+lCiHsJCajXShK28gtWo1YLLBdMfUkZiSv2MdzTdbCQArWkwZwVi8Numu/bmxLR916
LlF66grpBQAsZEwe9Al2D2/36Oq+HXPEgwFQjlF665+ge1sbxrnQ9J468ruxZnhfI1/mnoVVEfnb
jLCjhBm1LVqjY04m6cTfxKXVfgVrxt+wMRjAulYSrDC/GhWX7cndabHUhzLAGN/4hVVu+i7f0DT4
Tjl/4f5Uv4ElOqBdOcaEyG6o14/yqmuHYaie8KcE1acWeMVvjvJ1EddnDtnhx61YscQB/IGa5J06
OnPa+PzfSxeFc72dpCp30WWr0wmlWrWYJp3JaazaDtsLtJX0VxbYS0iMumXmkL+5iMr8NUkdhFUd
tDus/23tnTg6LvHEApxDYYtx7OTmkt7qTnUCkuIaNGgu0mMRXnRfL55XucE/D0jWkvtQfkWR8vG7
N9n8rNxpzq8BWrahGgSpwOyQsy/2EJDEZXecApMbuSIIXcqdGAN2C9MAQMrqbLFozf0lej3ZUa8O
u/ckBslXrZxn0ILnxim2ldeOPnuV+D3dGWkoQkzik6PhtavqFqkKe+mdafd4lxxGRIWJx5KVWn0g
pg6rO3AwSXHiKj49FJ/8fRAvCpweELRIOoWENBvM7WK+W7l0TFQXTy8062EccdzpZfjogQkOsflc
dQbkcufx4jHJnShTCwv1/5NvfVEMbGdjHPzrFU/6oShK8eSN9RFYtxZfJnDsKNWr9pX8DOeBgqOZ
U5PkP1pgK1OneRpFNskHOARX6Ybreg7bSeUwUPIq/p5dD/0RfAWa+hpcoIlR3V2XsCHauou5waux
kzZDxYRo7GMYR2IbX+KFoax5zlDabBbTMqWn0wEg+EzdpgM2uPT2OFCg+jAhZ8TyROG87SSqckjJ
jFlHIKe0vxWJ46WKHenM8VAxWhPA9jcxhjYqnuDQ7r0/wmXn+L+Xc0UDMjd14ls34VqGbJvYrK+W
p7qcCzPsRIRUYhux/BRmUyZBTqwgJZoTAG31EPB0Cv8GX4jNlQaARm3H8ANpj2JM6SaSzYuL7tec
aDdNlAcS2uA+/HIGcJ/N457gDG85g3dVR0FBX86xER/XTWPpAO3fGuC1l4RCbAih3O0RO7RNGb7t
7TpsIfXjRu4Yt+M3848hTEBMXkRxvdnI8OyhcLSYtBbz3PdHXMLz5/4ka5540nf9i9MsYY88vuSc
pbqQ7GQe4OpMV3rGVre2DXMoEn9c33LND5ATRaAV2uHRw6FJa+FP2phsLz6lTZlHQUFgIjTCa/kt
+0cO9JmJgCa3CXsmt7EfYwmT9UWpVcu9T6CE575GPBxnTLxRbOdAy2FzmjiDIkOvrPAjHWg8UcAF
cgZbavD13wMBmFgpTV0Qj2kJMndhaxrNqDkazziU+0bGgqU2jrd1lxwPHiVzgE2GFsuh/2VN8cZ9
1UjY3D9lwazd51qJAtjpabrZT+y8QRg8KGpVeBRyqhKYiTcTZEEqoXc/gDQmcsqONSunvFgQWQZN
MQ8Nu91+qk6eybfsV467bIBRE2gpcI5BiG/ODb6NTCKm8YGGSIt7D38sjL95rNjmZSPFSlB8sKRm
CgQ9rp1Idsu4uSdeycIFbhTAcFkky2x9T6TLbkGdzbJJYjDrBW2XmLdB90MVxAhLXj8gz8T3uxPA
hb0hSxVHz84eHMLc2Bf6F0Rycsj8HjzZps3gzixR7rXlwfpK7g5OBdxWm1ce20/BeAyygW+tmFBh
FxHxGlfTUMB/txVKxy6LSCSJ07tIZ34sIRfZ/nPtiqJu2J3dqWgXyevZVz/NhfNjMNIlMhlhU2O6
+8otPanBAs5e1S4My0B83BZQDe4YvX0lrxUvWXEyaehLDMcrv55DdYrx8R6BsDEVqclmtaXU5oW2
jnjpHOCv50b+F0fbgBsctaCIPusHneDjWUbERIisLK7Zd1aFAaV8GaF7EikYMNAcJNEmn0LBd+N0
pHEDvwmPzjvJP5cotdGSk//PdZ7Q2NDGvlsabxI+DKl2GHqb11KkQn2+ns5UYHxxArMgq4w9XX6e
RgZK+I489RUt6sPAxADMf+cyXKsmrsfZ/aSBYfjcmpSk0XyXdACdyynZ4TS1KHtqHuG0uXDurOGb
buEOAwib7M2pLcvsNvS+qzWMdeM0yjvJc59wjwt9wuAhlnx2hH67KAOTBcC1A0HplazBHVv3x7xg
iHdTUtonhe164Zmc9tW9ent8D0dJTWCnyprAwr9qA1ZXePw6un0B2zfgL/MGRUpcLJrLJqn60Aqx
bc2Jh8fpFbO1JcJrsbmFZgzVymEJilUXc0JogCVmVX1UaCRXrMq5OT89/T2qtppZqAqntQiNJjN8
04rtZSnl+yjSbCjONm/NX7wRG67Lsj786Xgf0KbNJEWbFAJjVWY5NFXGfKi0GohpNB5gq6Pc0iyC
3w9pgQNd4SbHvhepVqEPeZqEx9d2/BYVxbeUKbtNaEZ6mj2QDzgv8zKmonbB/nf3evrqeZGT9RKh
U5wb1jiKm2+W6bUnzA8PeBFSeHS5Im0JaewiCZl5QyvEZ7a3JWY8vPeBAwPIlWRZDxKidVdJNQhB
VgJQOvFlMD/MahOwhZljfYmOVFTuZzK6GZdpKXgrrzngtOLNwMrM/OshJ8WeJtpyiDXF4VXWmMsm
WJwV8J3QMkAg2tG5JDCivzgEq9CY+J8NWr7EKi/TYqjEXkVxAbpdAYEP3Q6DDXbZQDiBuGLL1T5D
rgz1iP03JKCTNOyoCRiQ5NKWIXnrJmcNPXGZ4Xg7dsHJiGwGLS90AiJrB49r0IG2VF5TpcMkLTNt
I23wGHfDNn621GsrkDZCKIu8/kwTnCgBJLtLjfTqJSM6bdeTHoy3ukz2oxynfKumXWahtxKUboW6
Xg0g/v+XB7xMiFKFY/3wR/SQAX0dAudOYQu3oeor7bqzP6B7isWFNMNBbwre22RFp21uOc/gHUJN
5aGQOx4P/REK1imFDN/kX3wON5lYyNn95lQ2mE+JC6w2FQOeNvu+totY/he34+6Phc7zXEBs6bNa
4J3YA8ZFHQ6OAR3aNM5vN2GVQ0Sm7GgBkBKP+TaqI6MxeGNaAOEHR3sHFnL9WXaHRMEOo6hI1+jg
CuH2Mw6ZxZJV7rakY5oo4h7vYawXX/zIFi1PHWgyaK8rycfgin8+gqqSDgaAeCvCYlXMR2tYG1lG
B2pbo6l7IvbNQFsztHaGpn83HCCPFymcXK7QTeFkmMc233HhRLLUyrJBV9l0/Su5SElrqyuRHI+Y
fQGgHazimLjsI+7zcAiNmEnbkeA/JtpSZSAZSrtVQ1vgTJzO5jGdo5fKGftH+x7FlTZhJntwsI1J
WcDgUZoJmWVc1Ok6z1dMl2Alrnb0D3iBM2medvfpMVW1TfCxPYhuizcJ6Jvur5mMLUB2/K9s1xIc
SqVSC7OppoHkdAXWTwT5WZ0r0L8BLTgID/CipfVsOF7jfraTrHGt9B/Ox5ufZCc3c6ZtgdAwut1N
m3O++pbyCeiqRc1nroz25TUHdyuxkwpj7PNQk2ZyXyEzP0YTctx/Kf1XbWx7Aeq5rNeHo3aoS9Wr
mjRmuLWl7vL/gds+x6gBWGaMRsDW+AeYdQNa9VdCeiBjIoM3VBQn5k88DqBGKAI0MVLt4SIKcAL6
YCjwTMA49BLJv9OHhq27G54i1H07FjylhkVQnaXsiz1ngJ8az5fw/XJ+T5OZKjHCkh6KsyoxhlGW
Dx1qJnBwmu1/G1hlif5zsXB0a0Esve/mGE7JHIjLMslmKXOxZQpbN+O1wJXDwBq0Rj5NqbGQ5c9g
2Z7srQYRSdTdIPxYLLgw2jc3yU/GREPM9l1hmyiY0qrZSpXToFFGE6SoIDYAk9NOFZYGYJRT9qsg
96hDCK4bDFbo1XVQWbuMoRpaY8vTW4cQXdUTC2HNX3NYmrirwZh/8TZfyVob0xVyIfJUTFHgGgVM
sadq3y5nkK4e0u0IGkkTCJkQJ7nAtx0s4PSzi7nC7ochCySwFkJilBvdULXY4FmG4c3okZXKJ7/+
vwVQ/GJuwSRtW3jXk6S62X7m32b9BtlbVsu+bsIjqSK5uAto9yaTJVYLONw9A4gapBLHIomtLEmu
ohzHIr8sBt2pOvjfyiVzxO1w8uqxM4Ko7kyzAE2hwbgnzORuoCBbDt9VBalWg5YhTpwW0aOvIE0u
4vn+9t9njtQv6EJzZYmmy4g4wZQIY8HbX50+3CWTsmrGYEfssvwnm38rINPrWCdQQvMMvsNU2vff
2gBNYeQReIgMd/NpiDAmiDRMjGNtwVWh0AYkBHQKxOx0xYRN5VdiQEcbE0GLkTGVfUjc81BodHQI
+Lpo1A4K78vYGoxrI9auhmKwx5lyiBlGdkzSYEN1P+JwhsGEPNU5NceXpgTpfuzhM5/TkWKqPbVe
AK9Zj9ZKenf7Cd9SfwTtw+YmbylEs0suEn9zihx7EMKQVClFEDhpMFvIMn5Z6B/BqFDu+a2b8QtY
RosW4YhLmhIHihAAov9BdpxltujoKKMnac5soi/choCi2CX00pzggin0TPIzM/pvlfA7PS59Peb1
kQ+d0Sy3N90e+GfI4ooN5zajjYisaSrGLgWqIcuLMzM0V00eFxgMzJJaEnepPwDzRRUGW6cD/m9P
lHsHlKnzDuPRyy0+Mj/w3TBg1IQy4o86S+XTBLhKq1BorChLG0LYZD9Q2fLHxZjSuDEB2CmEQj63
RnTWO0OD8uIgXVrZ9A0Zsq00s21aqhvaOmdYJmQr3x2hswkOkhXXAfQ3a9uQ4umBKHQ/Y1EgzsAZ
yNdI6Wr8P9+VlahojzDkk0uejEKJok5tlgpJdA4VrTEWO48dMCFphjaYw6/uDrtc+ixLDKDfsgcC
9nSkV6gg7O/E62z8mb38kE9wic7JVUY/n3hLylGsfl2En+wFhjZmlo3/1FzTKUUjjXkJVS+uStdU
+rvgQIWE8296P7NaV4/04tu/C0TjKMqD4CJdTq2RHAJscPCoDjbMCiurlzwXdcgcXKt4vHxhZj96
VGYpZxq7vFM1wVJ3EiqDcl0nWZqoBynBHf+dQ9/S2MDIoSVPxUTaIHGLHWE99I/qcxiNslsMRha9
2tw47D2Z5tlS9EpENC3G1+JYQdbKCnRYhhHCJuLclqsvq4yICxaNMrlFvcmIcAExWCzcnD74k6Os
7d9SFOka3P1Ehhs9TcbxOX0weN1wnCtJvBJqm7fYUBf/MNtqeoZPkpEhMU+7p3vy3Rp8epGKgTw6
e5wc8J4IPujf9dfvCKS3LZk0dQjsHk3SeiQWrfThqu1TP6fzo1d9K+MYYgbnjDMWn+gvdww9B0FS
SVI5n2FkB3UegzGok73E+XN4JiGcqJMSMjvrU8lHw737SWpxygv1rJ8vJ5TM4oo+r2T+U6hylceA
C9FFg+Ls6gyVIxjCwwWAqrWLn4bGVYPUrQ1c9aTdQKE6+tWC5eGKTknJrr6oOaiYFEMjDiTAk61m
Hcr+Dcj29qTVqnjRDaE0kh/SUMxTy3JG5H0BgIcbBT/qHoHgsVUd/O9nMkbKYGVVaik9QC76hzya
v6Wa5ZNkRSKAMLxWcdcEGFXt/ieRZbzZrO+T1Uo9id966Tkjs0P7PHE3CblCql+C2eE+/1Rr2idI
pPAZnwk//+42eTC/IqOe7JT/+AwXaMyKLDaNjlPWZGcWPfcR2khGTDFmRbCahOUxQ6xkLz/xjQuz
4Ez1xvmVpoGiW28AaR6+UVxuD1+CdbX1rU8c7MSZfX/ke0H8rxJdgYVHC1XSh9ItQVEOfTtZHwxL
xfp4xTk20gYoavrTq6t5C9fnJ5mcvecpIp23/jhZzRijJ+OjE6+1oprXNs2WDmnj/tF5biv/Am7S
hJ9rCtl2as0WXBIFTNFigOrgQPksmufdwpAPRDh4EvSjFu7BR/cm3RyavGdgF8RiBifcGp1/F0Ld
PTeBMUk/iLEG6vyetcjVYXmlaGREz15TSKcAbzbZtWydyoXvZsMGNiIuPmWIwptMgqHiPv3myCMt
ZRzvm7C8YA4mfGrGUSRKl3XEPbPlXjxG2jbHWNvu9qOYLRfLwwtYbFyLp1XZ1Of3zrn8aF67xezC
JhzRbBGkJ2frtTUkn67yY0Yu1yGk8zCpIJlycDZAR6K8+YOeN8MmeIa0vRfI/8wK31DRchySTOsa
yarkQtdlqClXQnxvPPnAyPQhQW4NlPt9WWNzq9zFkacWsbJTq6p3EoTXbyPeWfaK67xxqlOkMVPK
pF7NdCQ3GRab793D5hHZxy786sX1J81LdPeKNpB62yv6dPtNsmt+RoeHMenHkGWC2aSCN+zoSIWQ
nsYgDq9SUixfWCTg0JrUyozrgYILHsgKHOR+RbQMtO8eScAvMG5GGfc3eWP/lgxLpKP2PzcBZqF3
zVKz+p/3ANjBOAR9Sc3Oq5iwbM1E/41Or8AiJ3wKw59y3Yhf4O6RzaxxqAhuMNq1gKbOxnzzBUcs
hL+RMsXR+3aA80eMeH/cc4qaUmjidhmOwe84XrHNk9Kmab1tD/v2i9Ak+4TCqP1pxNr2XmGXyMd3
heO2K/rpXdKYQUav2fJcjoUO/VqCVKh25/+/nSRtJtvW298pPCs19PLF8E6UHsa8V/yhGnsMAo7F
q8yqZznZs1Kr6/CFfiAX+y+zqoUHT4K1cUoH61l6lFgE+8kwlzQdUHYzxNPdsSPv1Ienjf9n5f64
doj1huhqFUWGgugpef9HZx9kh1njzzvmny2YjyYBL4/pkozxnD9/FJ+hDoyWAUgxKSGmsXR68nlv
0bVzUCyvslYH9t+BpPfcpFtLQg7dU9Iw20GPXBGkhMQAQGYPf9PuZfHa19413AAoSI8jb52sMCWy
ZrjftDLqQyiykHF1/TriclDN+QNTTwmrDUOW39/ncXybi5fRXxlx+jF0qq+kkqbdhkcD7oZ8C6Ma
WMuWEdaDdZ/RLyxB2+XphU0t8F5s743pCp3JRX1+76gi8grPDUPFYCa6jE1cmwCSyBddN6HQdyvs
LNXoCGRYzkR9NCwjXRXHxQlS8R5wsc80xy7UhK+gRtU01npjaHapzw9kYnFU5RmTBqS5R33z3k9/
108SeeYY6nIMD3ZE2baMhNXOS+JUH4EKNAFkkd7rhKQttPQCh/MNS73CNNf32eVl3tFZEAaVyQuo
6BFz6uvmsmuBjURcNEs+OdPu4EPcnx3tLUuhgpIg85ZIypCllzHByX5sqkwcfBi0Yj1W7UvUiQo3
/+r3AriuW9edQbrGvCgHpKWQLfGuWeOPmL+2qOh9zMeAk9d9Gj5mDaExmDpHX+saB94un39/gjCN
GtVGxlgU0KnbfdA23Bb037fBQyDe7iD59/2fEf6nAOV1yvt9uuDaNCVjEuS/Dy4XAys4cBdYDiQg
WS3RcaXpxWxOpUvem0+DU/VU2wZ7jmwK9OH+lpn+it+GXtFdLescInr7Memeu1BX738GmDQIyRt/
ZYQNUgZ7W+mPB/3xObWOkrnNjMTNw1+0Jf5g0d4ChPZyWd0xZ5Hq32P4++4sX+S9Y5lehYcKuNeN
pOhC9PmGp2gMwSXXW7VAQ/jWlEI35Nm5jDFh9ZN7hxzUdlfjcJ2KBbrMd8ebbd5HV68NuGfHKBLC
P1VTbLLGBtNafy4JHX5aL3f+zCoWGUdaz7jj3K6Ju5uVZ2IWJ7wabYRAmotUAMC81GE9ZclZ6+dU
awV9zrwZyzEwzCELHroJLvnamD8aFM0x9xQewlRHGYzHJHF1EL6RdgikeeZC+xPcWDG9aa5WWk7t
o8AdV0wqdLEouwXaHIbAYHRI2fGZuUg+fIjOYnOLXVeawNOklvsjTREa1z8p+0PJ/pCUC2vgySwW
QO3ILVziRqujgCAWt0hpZUv1zbQXUiSHWGANSgdkG8OCUKQYyLplT04IlqyoZPShhZ1HUYCI8yPq
5ZToz+bsEcg44ydkq8NXW+jYvZyFxBjbLuXrkQgPXo6UbzMspx5QEKFHL9yveX8MrYxw0wkaAnhm
KSxtrVPjjCs7Jb/bwXbVSVQKaUKx4NJ0GIy/H7DlM3pzywPFPGsqLkSAmSWAtAw6EQJUYWdPPECh
I4ar8qmhJJENffFmgu/EdyywMWoTnfmsuVac+nskh9joEk2etvcdaAQprcz2bIGDd8TEH5lvgl2A
pZeODZX99YJTnOi4JAwXLEfwzLvrhE2z6T4YY/aJhM1HiXWBT6L9VclafmH91jgIgRxOsxECe5F5
GTBwVL/HQoDBqtreIqVE7VEzmqsDGXuwYj5DSFy51L89AyJEbUrHmJxxkGgnynyA4pIlEa51zAAR
Q7NofxpvkrJCsWLF5BIpn/CsdjN3pXtKTRU4d/CpS3y/P2BCnW0bSOitVWJg9Lkb9l+88uloImD7
flw90HOGltGTnnhyfqjrzIay7JS3H7SHPhscVIKEy4ki/VYeI1H3yVWlIuCGQ8CAzBiDjBCc3ARI
Y8EfVSbTYC4WhYXaIXOSPEaNvx0gsK1vNs7ADREeh7jBnVigCnV38c8F+eQTvEERDyrLRAxDE8SK
QPddIWR4rgN2G9iRunhOl12RdpK6wKHw68ZVlapM1mwwKP23v7jm4ZhCTARJXgPcxywetyGD0KXW
rW5IW13EvlFg2QUm+GO4JzI7nNgILXV5PPoTuy3MqBnhuaLDmMbYfvZsWZLBqSNABC+mQ1aD41En
PXh7oHx+lAiuHESV8zX8NMB372C40sZK3qG0NupmDla01LRus0WQ2N7pZAEtMGueSJGGw3+0qkZO
JKXbkGfUjiClI5qWHUVExjFEnhAIyV4gw4k5e8U6NNBV/kY77c86Dbb6OTJ2LCLrSiXB5CXA5cA7
9PjvsqVuahAseeLblti5EKYDmPe0Weh4azd6LdGPp2+02DjMpBs6hlB6bKgjxpVZStMM+jbkSFtf
Jvi3Wf5pPVXejfuC2anyTlaYPYaON4wbX8kc3/ufANTIYWpL9WpA6VU6xqTSJy+6KBAqHRqPDrNf
ujAIh8M2PGwXi4KMO8xXZgKVftctWE5QR8R7qVzWgihmoVYgX6nKDJtCcnpP5QBZkEGaKyOd9H17
OnacqBaSR8yP1pl/tGcgg2VDVaQ4ELGJkJwET1pS/OzgY10ZxdvkidHxndJwmhstvXW+qbBzricv
d8QKbjx9ukTmDNPG6F+peNGE6ArMlo9fYwVa7R+iKe+aDwHjPQR+yFN8hI/U9iCOtRsZLl2X8spa
o0YevSLYIkt2ndVWux2llF6Xyq0HpPVR0LpiCKhptPhU2ORyRHlxtIgsWK2h9tZhNWMHYPIrVrQy
SJhNGH882FeznOzqT3FKkkIh0vZ8WZD3IlIlqKC4h8aTsI8AmZvllIEcVnCVIVpMFFJxjAgYPrrA
JeKr2RwLoYDdVf6Eu/c7cZO1j9I+B9IUSWbea1i5xZQ8eEGJYYF7wCTn4b2aJfGh5f2iRdAMk0jQ
zpV4hOaN+y+uuViYUaGoZPFOXZPcgz0yiWaZGjFCAsooqyauKNgknW36guRlxyQFMuJA8XdLePOp
SgTQfPiWIONoboj6ynYplKr3m5AcH68k/3oyGyGaVPjytiKRZiUBrvUyZocuvfHe9jqiS0zMqFCz
S+KH0FuMDoHlxJS4afS8R2EQv6MSJKakR8vosci845FWoyMdDjW3oMs/2eZLgpaOSPaQ705CIeL/
O/pgW4fL7Z/R2lgpyk0m7Kvm9CA69hiiZvV6DXJLy3MGErxCtWy6H8AIHWCuEgXvBZIu75TDS++w
/wlmuL6vXdy87gMGBgRtWekzRrsbWFazOJfyclQ3IA0ZNenNyoBe8QRk0gzxTkhrnKkhuqgji8QX
OvDFdAVRBeTOHQVIKQmcCmTj8SPyh6InL83s4Unl/HoZ0QW7uWrxMFR5rNnGfYdx2UP8AKqiq7KS
JLZvr+aepjLP0siWecAzmhp636pzbevlkpjVkfnTz1sHcqC3bJmwS7D9O9nzBqzT1rtXAVk4AhRu
RKbkpFKErB+biK/3kgrF981uhSBkjzqRsCoiZr9WTNpwiS41TTEejgmG3UUC6Yujsi0/hq2uNlBW
9GDjJ/hNEjY5re1PHVjRZGf4qD9Y/JFavpSkVcNAa9MkSDklll2pdeeh+hovRZ4IijUVEyMi09bg
yH5yivdOx83m4N+AwaHOEbx4SVVqkHPaDMto+h5DRZ6MoukcgjmrGT/lTelMsyzXayY0KyEmfGr7
RkMvKlgpdCzOb5gVpHLXi/YyK4AkyrPOCY609ZovEcSdWWN+o0oxP9SoVoaeC8TpUmxSu3hQvL5s
uyWqFWtdnUNEqwNdUACgmfXxcM1OHGZhuNa4g2ozsjoHOAzx8hk70e6VhyR7/k4d+idvdzf4yD9h
1L3vvL5BcKy3yJ7cBg33+4ObPs2zNtxw2RjOE0TSJ7bXfAbZroWrop5ls7vEfzl/9VjywkMn1KUr
xgVxezW1v7dYQ63iDms2fBnh5CbZYzUYY8W58zHN8LE3khe2Pigsrzx8OT7B31xhEIME6fLm6QDk
P6kD0yRMYASuT2GLHm5QNAA/GpFAKYrOGNnh/GiED9Wwnn/sI2HCBuMRxifl0DdHg2enJX86zoc8
6QIL+piEdJey828KtohSDeIsWxfQ9c7b7WXkq3gdym60RBD/dadNAwnjg7FU6PQrpgDBpxMpN8je
4SidEJwYlj3fQshvPjwMm98eKp4GLIk7UOqCADQMaDBJihBGsq5IK08ZvwNcEltqaOye/8k+3GE2
UcdO6NuJJ4rNjSOcNbVw1ckPH1VPElEwyyQ8G3TA503QeVG25Kzqe7e29+Cj8wmzxuShsTkc6/Js
bXNOxob16MDZtiBpRCIxFyXCKwegdUklu7JNadQ2z/7/XRD17QoCVoClFSu1DSgnzk9eLSLLCY56
teEH7hF7dvaGQxlqkT6b175BYuXqVGs3ghiKRLNRpaCYKQffd/h3u+xvFSNqbjF0AdKuG4b6cLAI
Of5R8WmZz7XzNyu00HoLq1u5WXgDHktpLF03JpTGouApBzTVwFlnKdAPG6PWS/zLmQZlg3kNtnlc
2kklApcfXE9sc+NZlPw9mDrcw3z8GDE5btRE5Jo3ApbGRmGBa6zBn8+LHK1cSnv2wZwsuuxU1ViT
HB9uwY/YQjqq/BUulNyZulc4FjWq3k3bkktrMym0FolwGq+7pCJhFutilEB2A7hMrQKUo+nydvOY
tLc4M18S4zdiLfzeUqf2pM2uEHNcJqbhGdhdYYK+RPQK/nfmDi21iBBHLWFKdd5Hy2eO4PeHAcyM
rzL5glrxS5d+sZR+cfZrWtMulbL8kaOgUaTy6xcJAFbbMzlPAcFFKTMMzt1Hp+dNYgs5jqLt9MDb
5wa0lPKSXvFEpYy16fxb79heW93EosyNFta9AzRxMkKCKnjcivt0oaMlLZKMK4T4KREJlfaBxlqE
U26mEnFx6yWTfCAslTCcO1bkoHpSe7OOgz1KBy6Sek6I4YlIjdl55tyDE0IIFx7aO2x5FwGZb11q
se44fVESIGzhvFrddPr8iowPkQpTSOHQBYtLUSVA78LYIOFDLSKD48ZWJjjrGCUoK6fnCtVMxNYj
RyaZtn2SoDI1Do5b/XqXyN9mAnU8gjq3ea3NYsXKyGGJWv4EaYz+ARdtj5I+b1c7VPk2TurokX7P
YNqWGNOYwY60qM2PhAedkFNm48RKJ60+UOKPQaDE+PUAeNhJzipoO4zi8hNfDyuEdPfyUVqlOgyO
dJgaHsMvQsO4rx+gPFJ4FfiMnIrhwAMPhAb3VOYLOMkbU98Vdjzggj/wouPBzulbNwiS7GBQlbmP
FWPVW+2L5WnAcBhhpFupgT1W++0aOQVEApkkvh6TCRp04joReDgXS+39fMvfDsBzs+eX11xaG4tD
hHd8/21Pts8iYMuJ8802/FhVASpzzS2UPaLLfUHXv4Zjo1DMUe8FNlprj5epfQpg8hvSnDAgF789
cZWzaNmd6UJ2FpCmUj5rW64V78VYCr7M7eKl8fZeD8z1F2lJplL472wx2O/iAxC0um9T4i58Je8H
ikzv4DdOYhjkmxFmXM7h0YCDmStBffAC7Cci8zB38wnGBNRaaFuDuDX4umgObaNwktgj7aDYE+Zv
Fekw/DYzBcTVYy2JgqhhztTpmN99w6iHgVqBzUFxtKyWegOZ3O6mRuBWwzPVDpWefjjeEs/OpBTK
G0Wu/5op4hJu0AlyYQ+1PGxEif+arScld79vU4woX8znlVVx6zPZhVSmfk0jHpOjkhf7QaD5Kmut
T1Pcwmo+21BDK6xdlH0a2woppyzO+iH1f6hTLXp6IhU/ZWKnFRYmxOIwS9SV0CBCqxOLc5yrP00J
j9Ud8FGKsbaH0BbEuURwH/1f2bbtuBjvFOErkCa69+uBBOemuNasA3jjjkj1kEV9bLcsULrGGSPQ
j7f3XA4TgtmPsZ/mRSet/c23Su0wyN57siY091jAHVTLbgDXun2MTeuOtmd4P2pOayDiI/oi3M0D
T0i7cicHeB1ezBNIuBOmCC+X2UoS9DZsud5KnXZ8iDtuaaxVzMBHP7nz8ZkwTJ9gWwJAyj2VfG4D
sXAE5CG3QS7pZ+2Wxh3+mOhCd9jFXqdt39BkH8SgaQOJZ/ragWbCV6AhYmDQyftCKbltTRzCJD1R
FDIBZUP1VIJVT3cR1ZWDvtFpOZEb1H3pcOtvGDQFdPLb1uMa42SfS0IuxqeA0WA86uJRFn0KUjZ2
bM87dcITSn7NqPC/FbihdmpZhjI3AF9pVbxdtR4U7uhOQXqkYeaP3m8rFRgHJQnK8pTmoSDNXGZT
KN9fXuyyeSnNExoPH7NIlBSVP4XdV/pEdjMfhjjntsNUF/DmzU8i/PAcRvXOg0nQYHXNlUH8b4Ay
CnFH+MZYWV2byVH0TNo+Fh04/rmLdT/w29FZH2zgwOCJbuUyFv+JjLahsCDthve/ZxCXg3zRVJSI
3DX5v4bA2hapwrvpHG4VYxLzU3NZzd307+CQBRs3eBMmGoisWNUehkbHkCFw2GmYy7580DdrPD8f
0VMSBwJy2/iXn9BcIZZHJSN2uTYT43PJBlpnm8rO4/gjaDCDuyh8jhwxIegqKmS/LbTpkmFuAW2e
W25FQA0URojLEq8W0cT698pH0FzocgOY97t4VPZAz6YwV3Lg1HJV12h6ctLcRLNOJDZV6UOMSf8g
J8w0TxNy7uRL5LdGjVr5VVVp9HqeFElAjsGH0iK0jaiXGZDpFQPmj5UK/Kacg3dOaPdAX5CrfLho
lH3pWtHIxCA9FQwjp8p6cvEBoLh9ZdrxosjxG2YGY3aDnoD649bjdR3ne8S8SqBWzFwNJ0yqTre1
G/YBjmBDY54/zCtkdablLbEbroaO/UPhJCYhjPgE0nI5Nd+cH+77KJsQuoUU+XgSVwG6CRJKJHX9
BRNH4rJsgtMBZyDfCrLuZewzKqnTKttSXLabV5eddynl3n+DIzmV19ZqiWICiNh4cKqAFPe7lL1A
ZNyn2S4ihQI9V+4ZWkoxK06GGOjaq+hZqGe+vT3edPfeygwhi9N0B+mHY0xXompQdP4Bjdc/tbvV
es5LfHoXkU+FDz2xOmFR7cxpLufzMeI1uDqRlLWRoC7S+mMEwHfnRuNET8pLyz7NcA3VpyHZVUZS
+cuDJvCoUlvPSxoLOUM7U8Ji3/lOOMmwWa4PLg2iG5nlcfVpn70GSerIkGSi44HnHnWN3TiIMsbE
BWEdNx1UnzMjfkrm67DPatcJwtMZ4u/E4/G3gZyJPoR18rqZKz8PjaOvVWhDwPgl6Wg8ZDeUeU7r
IorOtEwQLBmyVvEtRyPG0BiwuBGezitSfQDM0LB1IiRkZ5NZc2kWmP0L/ZctIxcFVHG7xLmTdOk/
0kSngjv5FI4Y9+L9fqnOLtSWKvSWZazhGH0thtIVyPam9+dwPjNqqY9cgXMLir0u5CA0Sbs263qp
4AqHf3XHWvK+UfUTCF5Yz/al330LasUZFCDLcZNYhxGlWk2uUQEFUV5pJRa1SZd24fcSo+yQbaFU
Rnka2BLwWxrKWsqno2zTMCM37lvVJlFpVSnkjT4uGiGPtnysmp2TnxDnJ8fZH22MbwOrebryTd9V
TG0koeSfkKrziBIyFNsvLYlNC7S2+rDdvc41ZuQKIURibpnkJqY+WgGiJ/m79ZZGnwKlZD09ZiXf
I4f6YGEzh9CsVdnHdiTdIPZFKtri6b9Jcs7/wd4xL65TA3NQ13p/TuCSRnMWV/AzafJD9ABtvtuf
Zth32Gfj01lpD2Azo+eMv7FJBmfnuNAa0kqT7snXIGyJhYQmA0xZNInRBSiqcSgoDy+jK4ulbtWa
n6VH/2A/w3X3iqehQaX0tZcUZ6j7GaqtPzut48Q/cXQ5RM48OjvNNYK9w8fAva9gdFZrXwBmi71B
StHaa6lHRXjrhQgxAAn07EFVb4i5Fs5ClErxSmgbgSM8QBqYHjc+ZeuG1wBKxlrXloPRx8+DXWuV
vTAf0rW1notLf9odl8jFCDHeEOQU5QXDLTfEOw1uNlBJzrxtJPPTAUV2U802ixj2Ozmf39Pexyx8
zoK1O3HCp5RS7h6Nvy5rHhs6Z26bHxYuQu94H/Syfn6Vhgdf5pcoJyr7vPSSFRP53GOJXcXv2Ttf
IY/efcbNKZfUbtHplW0Zu+b2JsC7QQLovw6mq/Ykqf54tzUkf+uGj+6W+nPjDVizyvORIYTXZZB9
eeenP0jr3nt23QY04h2vAQNpB93CtMUaagIkGXmDbI+CkQ0VPfLqrpcYvdfQDF3qaIKP3FWjaJ/q
OP9k9/WSZLuMbAFWd8oA8+4bwV9zAqeWjgO6lHbrbw3K3jyP3vlwrHP8LJxzVPyO2vZ6kfJSQbgC
1PWAMaBBMZNuxihwxmlhs3gZnSENiLurRDVCyuDqTePLeakG3nZDWb6F86hIK5JaPmQAH6/2fCad
2MYes627qAS4e8syfTVPAc+htztQZCNHY0/3sPJIphww07oXhUhIN0WrX5oq6DRc9MaCjHmy/MAs
NTgntmB0tGNjUu66MXyUkSaRkbv9wMmHAWE9aC6726pyePcT7QtKXQID8C/oa1Uikcvb0fN/vpbI
E7lem4N+DcPt2RGmwt+tANy/hEHpdM7LhyjCYkTVq7RdzX8mUsuJXeylqjBxV+GdXsyNnkl7ymOo
wRR1flKMvJaFvnpBk+zoBcY9X1PKYN8z8qsE+3GQyPvQ5YGYyEPyys2Vo6tObab4TFpkYMlKR9b9
0hKKV2n43x4k5PBLL9djvTUAF85NZlA/Ax0qXEbNnVpkj4yzWUNGWDgXLJoS+bf53f31ttaF49KM
7aVaYfmbxiRqG74j+d4wS6Z/HdPPdTZxXfiLtx/pCdHwnQs6lqNAsB7TGjJULwZGY7O+MYTMP7Pl
b/1ObfkuV0MOC0u+3MxZ8o785/U1AwhJQErPFMI+nF7bsZdmX6cG5bJ+EXO5VyIgWIQyAccBrfz1
x+slXMirTSZMdmyIvVfbIC5x2Fr7oBGqp1fMLqtWWrBF+G3lizp9dV96pBzwp/vb429nuZ9amxN6
WP83L67cWCCLhSr2viqaRfgBdPFoDQWj+qfLOEaHuVpryltEzXVXHcq05s6Ihu8QhUGDKKT7qAc3
BgWuHR/AVSbyz9bga6idkIZ4bQYkI4mHzfmYBl267gs1qJL3Vl9jFKicu4L0pFJ9esnD78Ikw3GC
7j4G99RMQznSpChfDF/P/XYrNdgdVd3syreqxNV1VIXSbsVcEA6kLTlwv3MYWLN9SV7TH8/eeITC
lY/q0bR+CF9cx2cIjskSuaBfD787vpPibdKcwfBe8oJibakQiHqUDzQm4Q/K6sEv+4ogtwq9+HXW
el7h38G/DCqUnn/jPPVEBwZ6vT0z7AjqckyX/vizmVDSbgRNJkhwL7GNNRmENsWt2KJGaja16WYO
dFeMsG9EMVbKet2tNyS0h6A+1OddolyMpCJxehYpZuG+0wA1509gwbWKK/nhpgq/sEHhRyZN0PhG
neeoNh8+XtJ8WfwLgPQqZsDEVwhy/M1xsu08skIqb382hoclNo4kV6DJpvjtCWOA8bcFNTW2icTG
W+3NQy9B93oeaJYOUYCL1yWPmVPFSS2Fh0ld94Y7dIxu1ITR3IDnGi50VzGBUWNqZZ9DB9T6kMY/
CVEnKibpPqK9EXBVuyJkyKmQARqyaYM6QF0DFCfYQFR/KEt53/IclPOMa1FKBFqSQvKT4oUTHG/+
WNudtCb0y+dkT5QjH9G3JGhJ8beVb/zhz/hyd5d2n5hbSque8QE5v/U4uamCcwqLqRSOaAkFuUAr
OiNrecOCx0RhgX3XSML/FxysDwKrqYNSxbAHYLQxJT1Z5hSe61ZZdCX1H+Ho8wMUN+B/81IKlgt0
Ik9Fwq7R97PgTFvG9ftFAIWp+O73wymsHAWXdA3EDMx1lmwy54uUCMlCmhOrbpgdlzo034Mb5cLb
Ty/77bs/flqMHquMoDxG2t/ML+f9HfCUsgi7T6IR/tLdkUg5T52x7Nhj3G9+iQg4wOjV/w9B/9Wc
cvnFqSWcKFQQzDW7OMZhHYs0+HedJ3mdTWSpa3dhsX3rpYOV+pCfXhNZ5O0vwZH80hBsb8p9p/7x
HhnOi5zrvyDLj5hgNS3MHzuE7mK28PPhGfqPhUEBZ+I88V7e+PdyYV5v+r+q6zh0GOHlKLD9RRVG
fn/mTxe/YcZEjepjBKnHW3zlGBLij7iGqTV9IT5jMzkV1gUf0Ancqa1VxvGsdXUtxYFJSGQiie7L
k3onCnhXO8LUfbwcWlgRd/KT9Cn6k+G9kdJp/FiwI2+MV5nDN4fC5tIoS6Mc1KLllAaWihFm07sF
3Aa6O7HhakWtBfgm/tI/RDB7HwT/qyVEmd7BHIcjk7iGKzDCK/ugBFFgpVHWV0ka1Jtp5riXPPbh
1b3ERN/iv3MdBf9ddtXopNAwDlfZ3rlU4/N2m70zahKFIkP9OO9AApMB41tcrSTPXwzBve8GFZf6
Ezymd4CVRHe2gDIsl/ieKE+ZWhf5O5946S4Vn+NltY9bepxXwUm3Oz99V7a9Dxu3HCo9hoePFgXC
/DT3y/3u3dqJ+cPGafAh4CCfX5REjxGHCOUDv29uPFUfQ+L0BMBZYLQw9lGDJKXZOdAgz0OMALvm
m5grAWmkEM03Foi6OatD+IJWiOmY7pdGIFJVOHA75Trqzg59U1AqgYPwIb4xJDDr+tgImaScJKbE
9sH6sw0mfMSXWjoFc6UZwEwH9LcVxGwuIaMLrybp1KQ8nyPSOQStpVJj46erGmQsyhs18qWy8DTL
lczGRp+NWvqDn6LQ0q77psyWi/rttpWpE0E5ND+h/R1h7MxTcxGGgyEdS26ndZZTACeG+BwSgfN8
VxV7jdTnwHSqjDuZeCwhiL5zsiLTViO67lkxpNRTJIrHKfp8s2ePIl+mI8qcFDP3wdBob93X3Xh7
pdtDGkDA2+ExdmpfvqVhp/f4M8PDB2RmvdHnMFg5VrHM9kkSWa5gtP3Zvcpn5Ei/+JabP9RXtVVL
L8kBJ6nDmIDHtGfdUD+j2zu4voEg9krUugFmiItmuyH3QHt5P1+Cp+xNAYCHYci1UClTNWOPJo8w
OK/gM0RTbZPw7hzkKYzq0LvDmiQnsOIUYm53r33BkoVcCBXPlstYC39bAzCcvM9cotnOSNcs+Msa
cTT4GkDcYiBDzUY7q3gVOt1EBhWaS4+d6d3itgcARFclFFcYAApF1GzQ9i7+97D2YHJsdyOnnJHG
h4b3nAS6GDkUEN0F937vFWZwuhdeu/xlMUKbSk60FFgHcWtx6maOg8MYuEOsvZRTffTt0PeUigt7
PZKoqpCMDt3YAbLtxY2pla71HA4+hMQQeDd8gX9mcYKo/lxYNeHVS5u/p1ed5T/d4geQpA7uOND+
ZUP70QmvZKlHKTu7BE1GH5acIlEsY9xtz4LAOpjUVn9GEkaIjdSv2Ys+8vx/BEPVHi9iFFjiWqwO
1w60Zm9iowmsc/f4UUEf2hFoJ+I60FDXe3CCwXTzwW/5pMR/gSJDFneHlpc5abx0nG1W/hVx6iO5
d8wFDaDbMSEc81r3QiwB69r4Kdno5++Xnyi8625UKyA9dhcVu5SDGwZdsv7iWMkLbMzSDldm0PQX
XguKbsy20LDe0eeKAfEPaVvC3Op82gTt9srClFI+KjPRTGS8zFZZcmmkCaSvhK1N5RQnwki1ai63
58s99CiP50w5Ch00VcauzbZzdEiAwn2XzwbyyZbx+Phel16FJhdHeZCTNf825yN8KatZYaJGh2Ki
UrAPLHlFiUhGjUBWJOnzTqauOrnTZZYCzyaZIWaguJCP0FFHzrUvN3WiuxbtH9WvtWJGJQ9tfpfA
7LEXAr/Ow+E1q6yWnMFiZMIno/snqR0eZ9+fUD1tYYwSPhPEF1H4TqCUIUF7oHu6G5uCPBS495VH
8QDjY2TZAR7XkUjiI92ed7VhRiEYKF2QsTnf7ZhANPyHf785Pe0Xirql5+nh1IIrCfwKv14SfTzt
YSLsDapLg4emyYmI24j7OiRV2R1gjLU/0vNtQCXXQ7AYtEhbRxCggzP/qzJBmn/n0A2m5Io95L7i
j4FZeytRnFaeHBcIpczFWpgQAHvb808LVYl+HHJN0SsI/uIkLSjKCqOV01OIFibdNnD44bO3y1kK
HCcda0He/zM5OFMpb1kLl2Q6/U/PilZYDXEngNBxqStO8/r94///2iRxXYZtlU2uezPJecjelAs7
+blbN4LxLSdhdaJTckQ88DIa7b6PhiVT8D02dxt5r0P0CBdMdNk3oeejcVqFCK/y7nVD4G8f5RIO
M+Ks9e5N4RiQOVd64eSHFVt5rMuu/mhJ/7APP1yQkG+w1Pt6M9kzy/n7QTdA5S/6dX/Mg+q1RbLN
yAIDST01BQczWWYMwYR/h4CxHoV5BvGX+29EMRIcnmSjozTVwmgo1+8VyshLqvomwPqkinZOP8Pw
K0zpudDhy7L539R8QmNu/3dthvTD+TZWhlcDRDqtYzfWf4lyfuhuPe+bxbtjuotyuNjPrEXLClCl
MzP5VcbFlNKOtSu1qcdIT1dRemnz8KBXyNGnYS/vmBlKVQFZuXLOMgPbN/OV+cTFBXV71VBuTkF6
ZBT/n3JMuO17TO6AkEA3XkE+dCkpke17cV1wGiOz+xaSKUXpnmHWGVBe9ZrEt+dtAtg3o/o1LZu4
kTw4cswAbkQcx1kp41BQzkxVNIIshGQjXn4cYRR7QT88Y5qM/xWuaGhKRcFWMS34AhpK9Cr1abxT
txxIz0pa6mkF107WKKvyOCsJ4vLH8MGhnPIsLXnpsDvNRYJQElMB5gAOTOUTUjdB+DGfdECsMDDW
wpCljytIhOAh566jcd53pCX9birnKCLBscZXMv2H5DyGjp00vz3YHJkqyX6+gEdOx++u5AxF8JZM
TLH15+WSMICHXSrgfj6+yi52tukhtUuFLeq1DdPjvdEJFRvH24fz0bCDG9o9f0+5UqkKGoNmMZVQ
2FX8LQ2zyoKvmSMBh27Zt4l7GDjfg8VyrbTnX98MXojOMzDhjUgmKbc1E/6Q5XaEjX3oydEQmn9v
t7MJEvxh7J0YHSDsPWW0aK9W6YHxz/TcgoTxE266vUEu/e1UMEv5waNZx4kMQs7eYq2ekkN2SrAv
xqa/J1shT0JXm8FK5WN8RFCe9yxY0j4zOYU5a2j4rn+FrcAD3bTx5IN/CKqBVWUIieDMM/77/jc5
WB2E16evshppWek3IquKIrJzpWvPz611zv8mwwl/5qhvQGTAJNTGWi1ZDHeyEP4lv1/7TwW88RlU
yDbfjZ8BdrgP040G7BCcqYrhOwmpBJSjRzo4vzKtBHYLW9clSeYyeYlojq47UEBoypTJDht8kl5Y
nY+5EsAL3YNTvVYFrDDXx+hkhPIHUF9EgcV66FAvERsKTvNvNlPogh07HTPPPYFWg3/i5kp0zlXK
hvnR92o6yaGjc2WFBEqUVDXNMQ8a+OF6DyjTNgSLZmew1kus2Rd2lXA1Bm5Kjune6MbHRYATbqDO
8owlHzsQDQPfUfeQjWu1arOQeDxLoYpeEFYBLve23IxiDdV8MM1nmr6rAZ62BlxpLJzIz5Ns+hHj
zWFZT0yyVxn8IjepkGRJyCpHsPsz/rjiCwYQOG0I4/IR2ays4eWTG95grty7R8KyXYVT3oZLB41s
MtfZq7hSoBALi4t1R3QpUSDXbHNhnfZQUCQpRpwMWdOg8PcDXSyO0HVVSi56fw5PVsF2yiiKg/7G
4lo24BqkOCcKCTgGrL0XZc7dMJh9j8zvzJjOtJ2c20AowIUphvObXr1TvR+jJ5lKGdgyaEd15e28
WWxzT+LD5EkrEwkrdf2Zekbot7z9cJDYFuF9tkYcIkBvzDCQNMttTsdt4jEeZRWH7qJLXXsI9hhY
9q1xU3bADPLTHPSios+hQe/tKSrEpHUGw05ou0SFGs5A3GL0yfnDaTeGawoZBpyCeiVrBLHwF1nX
cy7cz+tSGErY0UHTq8K8H6FM/weuypfpk2NqXL137nvqKhNbYGJTlYp6x4+ZcIfz+kB1myXLvNGe
CalDneX2jH5sEuL4bzWArvlmE7H26sxaPrWXN+XH4SI8tJqnLwWbJma2IVYoQ93N4CqCYXMlqGoR
qe85gFQ5xct4jg6nt6jNfgzQidpuh5g/hAyMjeJEZvkWKlEe/c7lw8C8tk/+5mgBfEKW+1xKqbtG
C/3ReRsGJNltaBYAWPIniID65JGacPdnIk8FR5VjBEssHvDKDkP/puJQNLLfCYEmQxPlXvsPfj4d
A/wMFbdkBNVEm30Md8c7LAhrA1iyQgds8PRMaQiuzjUE5m0bx+gDQZzVCMSYBdnXHM5jz0geAz4W
ncUoSkR31XgDqU17dvL0hiurb0ao6X2+KxdXlXAZV1/8IdUdOZl0Miw/tgU7aBH5P8TzobDkKi2N
6Pioh15HOHuYlKYBTX3kFnZe3DAsXHgm4uKZTxZjck4vO2iI9XkzXKJZDnMVZAnZoOBjAbBw3PxT
BZWBKMKJwVNKupaoo3hdlonkA3fwG5GbHWRZszAwGCL/yembHMDGkKdPF7b8bbp79nySoJHl01QP
Xa6bJ9tYvKlfvyek8Kdne4zjGqucE0YYrZ4Q2sCwVDFxFyUf4g3k+hhG+nWYClinNqD47oKw6ELt
QkxkzzibsnHWII7+R9BXi2R5IzMB9jEFLGfTAfgfXTgpoifoypmNMt/sSoJrBZuC3pDWMRbzuIxK
xRClX4UGpRmqujoyG0Bn1aQhs5KyTBoGlqpNpkfGS8MhjEOfShCSrzpH0kghj9oeqFEoVjdvPQov
wFSZj6+KoOl2dPIg2o0p0Ue1CciAofkxKBU0t4rBP4QB6K45arHPMaF3XtOWA5o6o2oi+XriiJ9/
eLnVLawwDFiV1S9VSd5U9QlNBfmlsSsFKOfa3JrBzOFiwBz0Fkev5zqIbMSDHxSfOiezWswZUw5+
uTxBxGHUu1LO/PwoTEA2yQp/66XC7ZDIIPPSJQa8DY1U451/fH324sMiPF1RzqYBLJFTr6zvjxPY
Ae87U3VwY5fGeZ7z3W59Xzzg4Xn+VRvTpaEujzm+C6DNTVZxOorrM8WeEJrOtSGhjze+LhsUvYaa
P9wFNSJL7X1UGyWcusy8nzzT3AQx7lmpa11sj6NW8Eu/KFfvYR3rOFuVdjG7cONN3PaiebRWpQ4u
GQ4q5CV3NBDDf5qamHEvIBgkvdMz2CYe5m4o0itT4FLg6Aa4dNdekOtUDe44sZFmyjMYgrXEkAx5
NLAH9INoxWg3U3GkNp4ZUUJQ2hOsOjoh2WEEqOUS5awH24vj/Ml3/00WzRmBVrd1Izb2n8ubx943
EuJBOpCFwZkQbTjchUD8v+QQcNxvYo2B4eU1qMxC1qfbthnnGNv3EdsAbSmciGvzTWm5fqJ/rVSd
WNavu0RcUl9ryzK+51UOkMCACVPXzaZh9/G6i060d41XPNh+hA8NdII1EPOu2I2S0IoEYwJHb+gf
VL/m3mg5gVdavEOwnoHL2QdqiQ8Hk4Qr6o9glmoDj8mZmQs1SMABcKvnR5+D6ud1l6JvRVyCj9nT
tsm+0SWEoBqRbU1BRY8E6NreMJK0cmgqQ6PVNRwicSyb/6oM1gMzmcUqIszMb3hd+m2QrtPrfrCz
6XlAl3Pfh+Trqq01gCSqheFe9PqlWn71gs/okfnkF2uAoSN3Mwrd1G2adc4M8Lt+JoqRSYrVa5bx
3KmEuv+crW3FR0r4hlPLXeKTisvYd/SOHaprOSTjxm8W+EjyuilAYo+VWAS8CZiZ8JcU5YJ2aq2/
gTKhdgoIifC1bxtCtBYDEJGwo2htusmJ0vOiwH8Br9AqVIAyfoXEKE70++Tl8IuGdUINDMguGseu
1EeOnMvG0O4K8wsTnwuttlwhLJNLViLH6hYRthV9fhAYR2fPWEyrsC7HKPK2BOCoaolarDURUe+e
mamVfNqNZ9h2yillwLD1NLJJkD/2ub8h9MRlDL+NdGFy7vdY9JbUlaTbW87i2b+eMdNH6NBoAREh
+9kRRXy7K8Oo+7m5MEW1yNoPTuw29av8vy2Stz3xnrubjg4YWa8X2H8NniSUh4FRD8cPzlgd4Y+7
bITAkGepq130xNZDhLBTb2CVeVRYARYpxRkdsNaqO95+RIh7BeaGd2tbsoH3uKbltfDX09tbcT9m
Oa54iy/C4SqYM+0Lhs9+L0vk3l8Wn2oecjbt9beKAaKhHN+VdRJfEZ1CA05ZxIG+qepeU22DWBtt
XAlN6bFpp03i8xYJ1+S9fpOiQNoULNdoOkEFylaWQnGTPNKUhxlASWPBTKEb9nKLcUDGi+nrMADC
nMQ+ey5mmIvZJtPTzltcy/GCCjaoCaCzmS7A42e4PjImPyr5Fz9sIHunXP/C08AJDu42yqaZSB8K
lYwSJmVFIo4Zx8zEbFkRZAdq8bL+stpLq6+0ZSQCVJG2dyxvPndKlIqZDH8UUU8HQJLKPkR8etMn
7zM3/7nOMfOu2q+1DFWRILEvq6VsNkh0ZFRm1zNECFyEAn1cPVzdbesQe1kXw7Ft0bF6fa0DB34f
pW4KcfaShZqr/TracUW+xseGfkwCmCpWbFqMJnfBiZtKRoZVrLvpT+pSNdcbQI8tpoqWnlnWasjk
yqWDoTkIMckpyUVbdoQ0o2/nLY4PvZ6thLaVdEPbsQLLS7mkyv54fRBGjqUxa463tZ1bMbQGEqc/
0dv1lZyIE6pjW30UC2RepWRgbDR7ptH5lWvhtxm4lB6aWUfOvRag4IvkAEdRocfRD7W88L2EEacj
ZKqyS6S3/l0efXQsnA/8x8/rU5LHVpxjOhJ80aMbCHrxXqH0q67dtfHzPHkQfQO5jx1FoPn2jn8E
nA1jjSyaHtLdkG7o6q1YfRgfS3ehv4PE4nRm6YP143pBYkwB1tBznLewGHjcPTHWHoQ7bW0DiPk1
9NWTVNKJpgGn5Wz5aLpvwttmRs9xGXses8s5/Fmt4f8w4gowJFCI8YHmvMntrdMU84jP9Q2N6+E8
VSG2/Uvq1MezcpsZ04PcjfgnfGVt5z23Ud1YDTFUQaalaGHWev9xgELPr4XubNIB7UsN5ktjuRdc
sZqDzkXS5HpLx0QbCwJUO226bGQdRdFnsdJXLIKAzn+Wy/Eb8947GNTq+47pZa19uFUyQHJNCH8D
YErY900p7E+ZM3haVQKu1LRsrKvkJW+6YYsaCH9oIl7QXbRDdNPR4P28FIvvnJ8pLUIx6aoEI3pZ
pNXG57O4bYimQl2TW3YpWb09/MvZEOmi6AqYBFt7rNM25xRxyWOhAoth1PXFfZ6wqtTk/GG6kuvU
eCahPEiaCwSJ3biW15lP93YuxHilI/xwjP8S6iYvi2v57jCKLQ0CI+hO55RkQegwBl1X4HfE01r/
HItFazDOHWb5UIAT2CIFRFk0uV+kd8G0BIgavJEv2WJ0uuaKEDyGUVok52Jl4lSpKYasIVpDKd+E
FJwzdI7YlHw1mjCibFe8oIpibTbscp+34kVmiNVRBws337AYaH9Jq7AxwYmYx4T+PD1jjU3spMfQ
Ly+njZCx4pA7nmpDA2f2KNTE7znXhhFzWkQkXuEgR/rMuBx2n+xKBM+Rasusak1TIGBqwrbFYAjz
KgGENEBI5bAXnTAUE5YCsWuiKZn+ALZNBb01mlBvuV0hRA+a53tOGm3BgpzlqUzv7FUA76edn49u
8w/U0AQ4+xDJ0li5QuVPiyyiiJLhe9v0AP4gIT8VQFj+L0gxrlz+m0PCSlnkPIjlUKP464XOd57A
FUUU87YYBHbwd5UZYoj+nEbxe1HAy5g+JPFAf5PSLFbvR6nPwRpJMI1yIl3Qf+VoLbLCs3OWxGgs
teSKLmMwE9fQ64TKsv7J9NVBgDDFMVWSLvdSBoepuxI0b1MiIFy2vmSGylkHJFH1B7RhDJVqg99I
MKFohWC4aavxZkwJJUFxiKy95LmHMtN8mnBfjZAlqGjqzLuNElEOwpeqyjBnAMmtvn5FzKUqooC9
nMnMazNrCvb1JluQiAYafG3xGFfbBxFpDfO9ZAsoJOK4jlXrm0Pcj3brjL8iYJoxFu7zOPYbiwSQ
czK0AJtpyU1zkOIVhwUQD25Tm+fXWWc4dMe3LN/ytjHYBnP1a9Yzskz22OID6wFFk9hROC3l1zLa
8PKi478lntbAx0L+44QX3YF/sj3sfv5zqdhMYdebK5IM5yEzJ1UjE8mNbwHvKlMp8bz4XPNu851Q
rKZ/Niuue6ah/BK8Ox+aEN5eIbfvE/HbiAMUfLWiNRBr7Gi3DyW2LsyvGN1q7efeq5y7AM1jiw8D
MYpiCn6tRIwDaOeD69Yv1jrrFSN7Cf3HmDgHaXV4ytAwaoyJDmO0yA0xeutll3NVyzKKKtDtPj0o
cvcUUPIBafjClJ5bEfyjfheYF/GQwkwyiz6322sfenDbtpoQrkuHWOBFMf/Pr0wajjYxs71rji3J
8o1qPSCFNyiAKNCCJdtf/mHShLRbcUFMCsEL+r0DttMcWrc8pHCw1H9tR3VP8FheE9TbxxPsjIOq
xOSVVZoo8C8rBjQjlkKmNwsqWdQHytc+dz5hDy5iZjTo4Ey3k4+z05lwCIq9TbF//bmDSOres5Vk
daC4kvi4wxTQ77Lzx6OvimeqAzCksN7nHlIOERhczMev6bsiyfUVApins75qRuf4PHMhVzshOzwS
+ajBfHzviOw9GsEG5KFWic4RTi1sBrInuHqUzHQXJvSzXUU11vc/pvzD1dBR+ZSaX6PgT3NSD+q4
F3hbonuIXhw7AUYJ9lQr3pNCT5SRliZBuxrU3q0aqIUfyGXBMnp4ziTKWAaGlSOA4dmFhK8FLaw6
EUCc5pUonXIY+EsmfK0lFecXo8w4/jhV5FgKGqrAbpLENdfzZ+4VcGxNDlcb3idKwQ+1kM2iC495
kQmYn0mLwSdbA02pAVssSQ7p0552jmeuCQvEZdR59dbAYMxMpc552MKrYNUZGQT8uYSioHEoiKUv
D19HbKUEoCvi91sqGZk8OmAh7eih6ZYG06oaod6dmjtZFBFqVRChOgN9Io403wQ2mV6JLLcDR3YE
Y0JQk0RRY/YgATO27XDirz0apiCbAb1KJzIMjRxDNTz5YYf4lT55wqE86gSN1l52BsLb/xVD2a/C
cD68+rB2qtSLw5ap+EU8oms1AIywDTho0iy4g2GZ+QxHSVYROLE/1AJ4Hqc5JYsQ+9J9fzfqugcU
sichBqlrMlGAskqCMPRI5yTXxLsLjYv5CkXWknRoBF6xlK4l3LDfOT6q5Jy1wBtbq7qSevmOfMos
1daWpifa8aIEkTUYMr3I1MDeyluUDnHOprN3uOLrzVbR/Y+sJ41xg3AajKTh9yl6Ef/i4cT7lRVR
Jm+9CgZ2vdDcvx3y41MUPaqHBJMSvQYgl0yHipli8Akq7wEx24Zu5/dKJdQq5nBJ689m2oUp5Yr8
AzSbnwtXABFouCcqmdf8KC3a4ut0r6BBxWokggLTpw1m7RKGRR2AHNGuUUTP7JSFBvfNvpiUeoil
mYtKBTP8tEX3LPxXnFUecFo5dSK+ubyI44IdgX5UAXnOoVryJkoqJZSp1nr1C+zwiuUiKtKe/9Jc
oBJFotmHoVxsF1JvpdXpaXf9VWeCSvd+QORSu+/jBgVAMwMrAAbfh5oLJEnQGVnususWhzEylg7/
XPfP5Mh5pwLwjTuwASMqovtRaDIErr1uqriI+0bvcRVOuNf49oFL+7CzRzK4ZjGjVZAimIh7EiFL
DlVpSV0ag1yv+0r5w+ZV7TS6suFbn7HoqIpE62DtUzVN57AQBJSIPgMRcmbTPldxTulM1/C8G5Se
5Km1qGcPDLK6eAeaPG2T39AMoxwEEM2qDsWr0el0QhwlgKhV/8vbiS+s0jqwFNdBefKoNfoTmzNj
96nLJ5N0wH7P6DLsEVf0+0+IrD6ScIBwafTc4uc6ilkDiazBN4zL3FgnocjWkFO0LxjBbaFe1+DQ
HkMW5SME1z2htmSTe99CesVEkIwryBGg3+0NrPmvWXcbzMhwizGk+xSvDaL6koT8Zl9VsvwUKEu/
gDNqPsSSg/Caw7Lga7hpxwJJWlvyhizK+RujD8WkOYtUWhZ0Vm4/VYPTdXPbVD01VSwBDCcQoBJv
HCKtOfr1EFsfG/2A/JXn8KIqA7mo2GfZFdNZ3FMLgZlf8UU+OH7FPmTFJugg+0IxVMpQSNGV42Ec
OP8LeBLOdwJELUZ8C6Tnj25YnCTEcvTSDvdGHPQmbhE71u7v5naS8zqKbbtukV5CfuKTz+sb41UK
b+/AVKMxV6TDxqy0i5SLWgzxsh9VPNKIMtlRmTqvKAWM9IIOB6OWpL7aIk0aR+CNql01adJBOR5V
a2W6DcMqlNuQCC8mSfHXRX6Mdgxr6A6Mw1bEk9avzvUvbSwfArjEfdou6AypqByYGkZgdY7VeQqg
W4lJ4uVRdUQCdEsEhfsyzr4MLOENnvWucy/2Al3SgqVZVz6m4QAVa4vA/h8ZUyaQN+S+u5DzbRIk
s2nCBNE+GAbrpCXfqNaIrhhEd6ks1ltSqfNcxWZWrZuwXTySO35aX3K9v2igwZLU4iRzU3fz2QZm
swgdEprsrKgdrEJ7b5Ha7FfztNwiuTWtz13NjgJm5vUaJI0JFgJZCOIDs4WGl2ymzoM7CvkX8yTe
uA/zrd5qE9aoXHdPe9E4EfTEge7qF43z9ONGTF7+l7HA68LxkrZnTeYmJ5Ndb+VKqJBCrdbq6jS4
tjKMhhW9Yxa2Ig6PRKp+qtVY8VsTy55beUT9RI1KwOlU7tSj5HVDf03rFtc2f3T8TyY293u+Evug
DziW9XNegMPl970zLytHdi1vv2d1h0XfWBZU1umBemX+48t77zeBUADrW1E1ZVpE7WbWuC4Ncjrx
jxGbj591TEr3ZCpDewuSF3/xftIn0/lAclpqhvsJAVabbOt/q7bjYtvDw3W4DbbMI+hf4vq9VBAe
AKHau6kKrh+Ay8VBgvPCxYE9v4hAUWc8MzscyXBlcJwi7zFr+cQN+poRChiMyOoYhjq4IHFoByo7
yLerDFEBRjysQbi41Gt+QKUk2NIt9XR7qKNiMR3GsW6YQf1pMcERYtiylOCqwzurAs4Z7h3TnSW0
ZRAZuGIuYEFpZml8D20PA8zd13epiU35XsllnJ1QUJDyda5xKl/YBTTiivC6m5MCoGyyqf4C4vlY
ycaqX5eunlBkTkm/iYtKeF6KAIyoNl6fhdEOA1vmzZJC8+aMkBqlrxOfwQUL8cpr/7QUJAcH3Jfh
jBBvWo8m69avKduno7tMXLosaZcOXLkrJqEc3Ayk2MfiOfO+yeuzGTtL+1RU3N0CE8VFhoILZvpx
ZOhgDrKNVWf8KZhkzROsEKDMFYmnx+nbpitKND93UquSa4JZ0hE4FAQf8EzXi+4wcg/pnfVpgZ6O
JsYuJTeTHWKUZnOCdJf3VvH3l15T1QJDSEZYFWJOkTRdehB9W6dJpCNtrTCEK4s0yHilzCUCEe7r
ULeQExrPNkh8ZKzW33hwx2y6VZ+jmWLZ9iF8TWirMwH+19sfaALXfWVJR9+tIvq0k5M7u60maWV6
pN3HP34cqi96wtecXn5C/4teYOc0dtvDd9gs2MpcYX8pVZMx0iWvY8/qISD8QKiqix2Yz2NSYdLu
0MBxkyr13/59AhTNIA6OasnSf/yFA6QB1LdYSLPhmGQeV8v+J81kxWGvEU02GSQwBWGeE73CRq3c
5KPrYa6eFKgRKgp7SU5k6zWy2FL8gNnvUsCorlPWO7MFP4PobBi83kR/wMcY14xWdUeDoGXuSDgW
vNMltx9jwVcHbJzYJFudbjKJ17EmFN4NSkiE+EoaLBG8+EMZ3H8SUW/5FeHsjQBUIUqOlCzXepJj
o4ogtazbmvrPPMEoMd4ZDJCCDDC/ANHOyr4Y/4NJzFbANkbwcLmtZZ+Yk2n3RjC5y8IF3E5Il4tJ
tBfPF1QkTh4BcEYubbr0+B6KqVr1i5RYlqlBYi3/7BrX2yCz3LR9YV9NoIqSJgAQP9i9eEeJGI+h
eYWxThpLUmYO1CpoSfGRS/WIi0HMcmObibjMAJokXLEUmecW7xMfus3XG3i1xJ0iOvX27a4LxD55
gywOWLMT5KVnDhqc+DX9lSLBQijNsO2jNRuouoMprnyN28DkCb2+ejXJgSqU//B0iBTimM13YwOY
GtfX5fx7E2RB9+PxRb/XnpmubHFJiwt7S8+fwtqxkXf6Nr4YFG+5cWlEsL7kCHuxG5qzBJfVdhrg
8nt6Rcyn7CHB+DwEa2fi+Q8fvxCSIIGNcgUWUSFLHNwswLGiFSB/CffD/JTLND3BE5gl8yPh3pu+
AgJvvlT7crWCeRY3Dl2gfxHa5x+lRA9hK+SNUrHKBbKI+YWK3pvYN11Y/1kNjF3RmGPjN64TkULp
Jxv44wxuOUhtYNfs1nWyzlbNTlAkZgGxdUrJ6OsE2X9nMv5SzRCjFLD4OF1lcUGMRlwhSImnz0Ny
CKYSfsOhqqajuIhoPAKlWAY43p/RyjaJcx9A/tXFxF6j3kXXTN/XECqyp2LklDrXVEi9p5vAoTTf
O1iXnY6In+gFmC1gQSkOyh8UsCtP903ZcEpoWVRhFB76yvlG5gou1UBDMHYKNjHAs1zLWycmfi23
B8CGPEb0A5KMG/bJ0+jPjkwNBeiv6ca8WIucLBPXnkUwz06aQJz+X88wr6CHV+XwLPJhIIqmzfMv
OICAB/2FIdpJ4CtYnztu3JRlAzSFdqw0Q/J5DBbQvoipnUHffZWa0ORZy/KxndWuejLFob48mNlI
JfBM+n9U8vL708QVXWFHRwwYOngETZ+SsA1VsTvJiNrmYv+QJnCal8NJDeDDxcTCv2Po7qZotrfZ
dbbwdKfLl4/D3M/3B+ZbColONa1/uWJyQBNUwqUN+7TpKgwo+ymf2C9CUFh3asLrZhB/eELtu3lZ
oOJ9XIwFkm2BzOcZCt1fFheLsC9/i/k8uDMKC81n9vyKmldagfYCD6l0AxMK1YETVBhmUCq2VawK
czD6YpW6uo25v/dsRWFk7GcpGpI/H8aJB5z5tlvQfxa91sWXw/hTsKHMqgAq5mQZptfbHNY53Br7
ay1zQQ/JHwt1d8MKI6wTld2KsP8SWhVG9kC9I3uQAQFEymt2ydsVReWg1qTOPX7IsmG1QOMmQvRf
ZlG1hc2EWgdSRU+1DAg8xd+3qlxRLsAhlt/x0PtZa3/vKLBeA66n9kF8eHVb6c7AopNKGI8TKAGY
hoHUDOerffzfAIM85mxOdmjMLNXe2aW7z1vPsoqtblzmAj+xl5SQq9QmxSB5lnH4XIWcvL7jWrCn
cTQigsq0apzrAbx+eq/KcIwbS6OlV/dEHYjhs8kvtwGyfzVQ5HB2pbbSqYLFYW2UUI5AeYlPzQ9C
q1g//ABbuR8MFy7BvTAueI9xwNKGBQdprQVUxZ2HRuB2zoNtSDzNkmwyt340g1AUhzkKyZWcvESM
q1UEi1a90UOzuR4z7q/x5rZgzvjaWIQrUHBwguEtRdLG5KUXmrITy7whdMqoXqnfG1S/9dxRd426
nCMxFROmgdYnylljRtiOdHTtDFItv/ISry0Rt1DOMswRXHkeuMsIjTd7CfNLF4ClW23PdbOAqcfD
M40w0wKWnds7Agk9FumEH8UecaXJyqh1YMvNkscOw7Bd5MLWTjg4vMT1IdiMndJYYA/CsjxWgYtT
DCyEw71L8/vnVx/1dUej0P2LOpP3UTfulT10z68W7xMW6T+CaLrbnOtMRVxOd7Q/YUloA7m592fq
8RZVJJcVVi4XTcsJcZtNjkK41pBTelQd41269fKtLk7aBR45ommpHCrH4tH1ZkTGBcOcAEjHFiHN
nHVIthBQut/1Dck54+c/RU8KUMGflrcL+1ZnEEa+hky8Q0Tf4yC9SeKf1f4GxKd+IJqggwxcr6zM
w+wMfAwfDhajeXw0vpbvob1CY9/3+ioKWI0X433kQIRajP3QK/l3MvLyPyWORcdtuGhd6jJr1RA3
V6g7rfjcwCk2cMvPojrW61tfRJZwmRDZhb1bej2dUfBglF/Ovh0+s56sFglFUXYp1JEMUmebkBYi
XmYADoNYDOLZTW/j2BlhRrtkKwMF+aeiIAX0+MrQF9iHCztvzUkCCkaFZDs9kgl5O6BrQuL2HA5V
axzEmUaI7odBKGL+tefSgDM7PgC/4GhfQt8PhAhOvS3Z1x7JDcsGMzNWqY4jM0og4zZFDeUirpzt
THQrtp7IJhcirwjUFQEY67huM7sSi242pe5yHaJfvunKYezNcLUpGAJ5O2nuEU7T2UEjbl3Na2V2
eI8TbNp13VlU+iPgxib1olV1cd547yN1dCy89BgEuVclIO/be6a+XIn5h/sswNTR2uffmqmkk5tx
ICimVLJIX9lBVs3U5ZZE+xyYhoKjw/AZ5IsrMd6SeAwdD8XcoK/fXYw/8NF3sDluskIcgAPHT39k
DWFbCiQbZ0UTSl/ujR3jFSMP+v3Izh1j3LJhCqiPCQAh/sf0+hDzHGFjgmdqHQCAjTj/ujUhL28r
E0tCinjjOsmYxKGU2VB+wxFko1S7zb2DV3ZuZ3oMDEpXQWXKPbY4SrYjZTPZXoiw2TtwvZJoOm4O
eaTngnYIDDRJpqosdiKXUGyaL/5CBe0wQ0ICtP0RuiUcI714KV59GYk4LeuGiFVp1vpzBtnl87Nl
f6gmtwo5LvO7FFabeHa/5BeXwkJI41/uXx/5J2lWEZldAC9/lo36SxmahmUHv3Bi9jvZcfjIb9eh
rpRYKJm9fFZpbq8780wquH5m4oZaWvPKnGce9uEQOQLWahwTyVYUqXlRMFadL6pSPag/WKiG278I
Fp4SPn1DbCpHOU4y9pFnqnDBB3SxuzRVg2K3fQbXmauIRUtHrc3hh37lBAvrlxVyRQDd1PkcjK1z
D2z3wAYyAaceDjURBdzET0LX2zEhgzkJAGuQOKpaNgG/IxP5uDXOkMx9AsHyIxwoo6yIbr3p5wHy
jBB/KOtLLxgs9AyN2zMpEO/T6BXhw92gercWb0DXqa6GhJjpSp+NdgG2PyanWmG0SkmH9FvFnhOw
egQq5pEK6zvcRRQM5paqQzlQroGkygKyETaS8QakdzRg52YQ//1WoUa8WYGAinYxNk8byscDSpEh
C7OqkwDuXlBpzDcQNDD1pOGiParXD4bYe9FfS1ROTQ8IOb2JzbflOGntLuQ+Pv/C+EO4vJk74o3/
gyyiNADVh4amRvHo2BrLAzxOlm66Lu3C2wBvJE41ABam+TsgAmxd6ruCcQ/Wu67pgo/9v0pSrsk8
zyIwZ9f1oQ30DjzTQI26wp1KRowcLrBNgJP2f8To3zN05nhUfnPld74KK1xxtAND5xUK+r5ozT4Y
oQPHblm6x7B95OCx4oODINd2U8FZunv08VrR/uTekOawD/xUq5fixlUskQyrWXjCPo4P11PrICPA
8wKWiYIbxy0P/hbDBH5UoQp5rJhW9clc7KA3rIuw9mzfInE7d0zfVQEIsXIRoywQl1SggAYQ+Tsg
XsSig/zCComhtJ3n9HRrBlcHcG3s3rknIENgjkxAu+hGVwJ5UlQHyX0rzdwEVGGgzsH62ffVYE18
D79FmDMMzP7qrxfrgeQ9xyQr2Hg3bGcISt7513Ew25L1GAbDK2URM/xgGprflwth7f6nPKmbfcu7
ED5SWqhP0gvhiID9U5O0WImX060d7yD6JACBVMRoNBZ0C0qabVbdoglP7BQLBVF5HQ6DRmHtEBti
UrltdczjssUzSPrEsCqXxrcogZhMsIEG8VWEn39eueCehH1OelCLJdnkE3r0xqkzciayhaS2ocrK
Yo8H3pknPebf54eEkhWMlEm/OyKXB5CdxD7poqj80Av8PmGbD/jJeLU0idXlWDqyZgQw56NZKiFg
ZniXIped9AwN5Sk3SDwJs6IVv60/cq37dWG7U+XcPWMs9hAC5ckRjr5wUugERhadVlyvN9YyQ/T8
TE8TXNIUzMmZXXY+YdkEewGmglmOU3vkAOw+B5Wst76xPCRPHg9mFNunH2OpX0p/kZA/LDv0w72i
QGFYukzhu8SO6oGq/chB3ZeESAJbWD+Quw06Z5CcFID0/gyaLXPHelqLdNkblExQKOgxjNVzU/a4
KRQ1QHfYU/uO1ID2PwhAHBMlTyAF4/+ghdwWND/X6yUhI0xNMlEGhfoo0G3x2hSwkBfhgI/PEkf6
t/48yTX0BqxC5fHTf8aTkTw4GhEreQlfbb22hU4zuJXeH/FAISnpPTml9Iuxsql6efN6oTLNWXD3
eclNG5ByrolimVMP2lULfXAbb3ROFUMoofpfdLodZ54bjY2V9nOZivwF7l/oIieUD8vYoOtdh1jB
W5Ae+mx2pb8Aj1CK2tqSMn8jG0XVlUN+LJvLuqlHADDd/aXsob7VLyJ2yI7OiKHaeY9STeRjj1oI
jO4S3O/m0RiL6S9/qXhea4Z8C7CYvACj3ul1eOXZexH0V2J8o2BesRMnvQy81NLtpMCCXApWOTII
nAzwQ+GioM1udmfbCqgrv89ry5/O6qhvkH06zb/16bTnX9aPDpR2hwMKv3Q+GPMEszUAWiA0lXS4
tMt53mpH8huZVsP1vGj5xE7v1RmDk6ZsdJbmQtLR3fKGsz3YaeoNGS0kH0HCwRhhBLmS9uqNBagc
26+iyieEbm6qldj9ZuxgIWAO4ytGpvBYUwfU8tY/7BPw29Rg5IgLjgeZ14uPd+Q8cctkzIDE+5Rm
jXhT0E6MowphuCkG4hUNIh5PkdS4jU6AEKwJkw9z/Wqr3gQCalukmm+QfJwnGfdJeqWVNjxz6MDL
Fb4K68BWtLZgalr86uwRR8WR0SOv0WY76XyXkKVh019s6B5pooPnc/CktltwhM65FSAeUJSlDnuv
TJK+YtBqTXDs/JkxLxTv7t2ZyEpSZLGbI/afXcUjOl+tVFCgzhCEZbL2BzafB00jb0JbLlE6fup/
+Wixi6+VQpXUHohNHK5Xkro4Ddf6KimYOFnZN5APgGVAW+cP0DDGEBN395tRvDQMvI7wVlGDQYue
y5NAjVliTqYwRfmbJaeZHMJQnem6Uo/T9Sw87edbWLJB1X/BFV+ECh32bPJO74ynJ5+C3TWqk7Ml
P9F12Pm/s8eRHGVbvE9fWpZpSnyPwz6a+KU0ZyNYSWNx6edHLtKld3bAjUGPa0vEhunpJx36+o1T
qIWv9mIVUcX0Oug+O05ZfAHLsp8BeZsQygewFAxy0z6ttXzZuMcjslCrz+yRUdFsgZHmgM4vjvsK
BioxfRvoK+Yyz9ALVKBAM1Q8ZpzX/+FrnUBTE4JX0klfqsZm+daFhnO/CKKhWJypBO3jEJEG6dtF
t1EOjKwTBSKzIQb7LuqfFVcED/IHziCOZ4I13QkHK0ocgzDvdRKkn5PUdPfOFQ3OQ7y1vc+yEywB
zcpIfAGOWrjPtBPATPdckdPB3HzmX0J09SN1BfbEwCoPZJKRQ0LcdvHtGSBGV1+uAUTfMI9nt1Jd
f6qNFWqfwvYi1j9JpiVmciWv+1yO1vXHDTp2hhmyaHTCZB/jqXDbc8Zi9tUWua0EEkvVHaRV3RBA
S+sEw7vaGEhVlWnVVMAqr+rdXWndW3JIy0tMXrmCnKYTFg3eEKPSlcWKlqrvtSF00q4CEg0XCmzg
aRIG74F1DT8aY/njkS3Vmj1tO39slEgLTrV5c5QKKLmvonjpkqqZpfKgVauYdAqP2Q1cNGKfTpOW
+rJEnkIBPSOgyI7RUaF74IiqutgUlc7J/tWBZv9tk/6hVnmDrWzsHRlfKJ2ymfNN7Zo6TkoInWd2
I33VC5wP7cQGtaFWJgNk0yCmn7ZZkfmn4QhvlhBQ/PE0rr9XpNItcksp7ibS1a+rHquG1sUmAx27
Z5EIZ4DGORuYSKQos6WllSEzoc0gjStUrMLpmKJAGfLOIIPNeiwRrPJiqCQ24vrNpp5L6lNfNKCJ
U7eZCTOyKbRDtLiYbjEzBQrmHXadF69rTohTmZtN0JrzWCGZ0ORnXF9ZEmOFJ+14MQaBv1U6SJfK
iawb6GwfRJaZH5+Zxb9pxjiGKALxkVi+OkbJ8KbRpDDAHhIQJEiuab7/k2rXi3fe3Qt7OJ/qhBR1
IpH8UOX2j98LnA3XLiMiY7smEtbSS+Y5PnLuepHXrybv7LkG4S2i5c41Pd4JzoGbrf4+Abta3fx0
/ga7eqSRRUlKbL5teQWQTwK4kP71vYI+3tvBR8QbNASbOEraOqjyjDz68EG6SWul4WEKEvXD5/7h
uSOPJcIyj3GqGAgIhPOVGT70Akb0hIeBXrt7OLqD8wMIVLFT2iGuvpY7EeFGyKgyb0A6glYqwHxV
FpZLGlr9GRwWENSQI/sTgQAwy4/Cyd2iEw74X2s0fjcgJaWXaO+sGMLetFnAoLPLDrp9yTDFdaTw
80jM0fsG3ppWr+SZ76JprDFuPJA58hs6DKhc67IkKVAwv8SuNjYQ0y1tgl8LSXV9eDAWBhnQZFY0
TxbmGpwqDUNEiK9pZhwKVi7JlRlvOZOebee1HHGURbpy9ka48Da4EhWNPMFrSHYp9hFmq/6uJznO
F8FnNH52YyD8CweNBMzsUoafEyyy2zqINYi/gNaxi4NqjBywDiaD3/dcsQCBYjdKOHhvBSXqFfDv
oRwCAl/kSTgDLn1c/EGRfSgtAPwBOpo4mHhU8AqAF0TOHpvdFjEUq8lL3jVlX/3dPRgml00BS5Wn
EylSI4FkOxOAp8UYPt2sIHQDQe26EmZsJ0gpuDWzXhAlx6KoEiHw7EFctnw6Z0nEaFjn5po5yFEQ
Q47wJ1FveWmtX117Ei6S0iw2LjRrFywPvJoZ4qvvJTpuA1IBnQzzwMfguC7JdxRFXdJn5r6GGbGM
zOOo8Kmp5kgMiNL6ViUQiomoVfkkmrhbOzFDjAva4ZpWKNY4BSlkvlOo6TiTAph5RzWJD6PfskGr
FRqqBWB7hFEz0/MQ3Hg2splCiZI0L8E1Ap7dgXHPou9rkscljvLxTOu1qYhLGKSjbTnLru31N3li
Ze2qJgNXN/wfqiu/oPhknzs2+GAPsfMuCAzIMCas0xPQOi7tgfez1wB9I6W7ZbbK1qI7a++objyV
NugqP+ZwCIA+sksSSYq9g3RM6XQd/QBw2+jf/Ag5iOCT6BcZi12LrEKfIspk+zQeRLCuemUKlvM6
cP/hgrPh+4oZCcpQzc9yuq45+hI+lpp1g03ZRXKaMRfRNKG1K5qzRAkw3m30XIa520l99dBXTb/8
WSedA/c2lvS1CWKEKIwXJ5Shmf3/s9F0cnfbxwysuiYEgXc79N1juaogZbSW2yIxuLfy5R5lodom
0ua7g4QZBXG0lEAHrhYPD7OKPx5X41FRbMBGRCSZnxzdqWzn7WHgUR4oZlvsGeSHMrvf8CyWvnkc
v1xlTG/APCzMEx/YeBbMYaOe6mJ2nuF6NCukLW//2D1RB5bxknD9uIJSHDUvtX2sEUSeYa5jld5r
w3QQ+2cuE7IYcL2z8l8m8DzCl1XnB5zZHjq/GJ+2rdCLLYZ5GwFFf/fkH5GdPIooEDvuCOhXkGMX
Q9V5so8aZlN6hZgXQjTaxlk/9WsTnUNSZAGKOE93L5ho+53ds78KrJdMMM+EHswLywfyc+NU+DVa
WSQG7ZRZl4OUs7bfqCn3sLImZqXPV5tVttA58Rzg0Vi4KUHCslOai+j+qD5Y6p+p/K57hvCPlzB5
edIlk8/KWvxrp0LvTFGlorck5vbS3H5eU4ItHQsIiISkA/HOuKOUe/sQ/e58HYvHuKg8Insc4hVo
7C/n0JV6nfNSqyOdR4MFyYSiBUS4vhdHasOIY4cYpjdctVV4UzXdwXW5SVTzay084Y3hhkkpwwWA
CWAhYQStxFDd8AYbV0yaQGRZ4HGu0fWk1BAtC7Dw95ebLFx+sbaM+Cp7y/hMfRT/qivK7RvOOy46
1U5HglssR1UNeUn+AnEO2HZVt0hKmJnUK3Ekr34Y5sZ8eajMxBnWUz42GIWA1sKzFS91ejItqtqf
eMyJ9/1E97Az1JB9hzCI6W1NZMySgJOxwpRsC7pqhuRYEm0PFXimV3NVrh5LnIJCOhBl+lzu6sv4
VF+zX1mMkqS5aHtLaNNVdmIO3AbJxw43thmHrVxa8W5pRtS57eewLcU1kYVBP4+FjBF3s9E7uCmO
5KgWSGjoNZvcj6ei/dowV/4JrCZCzINao5WhCyVwypgG16dd201gcpODnb8I67g1tN+dHBRFxhg5
MSVJxFKo+nlQllHQxws6n4NCQ9gynNdvpfUtNlmKGp3gXXlrJ3XXDPPr6opXofD+WYxJR2DgYTcm
qae8L3Dc1rir9fIt73lhJiV5du3uiC3fqt5cttQxrXOViL7RvfuiFnC8MbJ/SiC4H2Nxl2PIq+em
XizisNTtW0BDowDXgw1A5+e2yTGNBda3rE7csBgZ1LVVS1QnNloHJf1XFwz9sxLkaWRhWvJ+Fjpt
KFjbDVXUfnxFDqNNahsQhDRLj2V9mq+YuHqUsvFZHoEyiv6EhgTDJaFPqILc1GgbVwH/YWKXXbPQ
hmknXM5FjPATyf5UE/8PCdkt/VXxrUGVolgQZOhQcECZ1JVNlwEE3zv4mqD2Gs24+gT4MBWcnjq+
Q008uPrdoyhuPBr1NuhS4v1Sn/PE9clUk1rv5oJsqI/sP4pt2V2MN/yICRNhn7ozsm43JTWJq8UP
8kEOihThG7FGD20flyHZgv+Y8OwUGjmIALBhZMF6JmMjLlHkhFD3H8i2fKWW7zgxv8ovtQSe+d7L
pwj+4+LnxP0O2IxdkJU7ydlPw+iQd3esU6dW0sFtToKjLq/sHEsQrO8EpwtCijPzZ2YLIgDuMju5
q5Nmsr7R1FJvYgQ2BiCbA+CBPMrqPrtInYU3zX5dW4ivt1Sp4vH1//Jo7WEYtzGsdGUIvij8o2d1
/EAHfPvdi7Co9Vzzkzmd0ukIU9tjwWbGk3wP1c87B06y8Py5sp0c/M2uV8Kp6T8G4Ms0rj8EzQIR
FrNKLqVUhrXg83KloBB1bUeclECqovYqCvRuvgVPZN/HFXZ+UJVxcbV058U75ujUDzEhkWO4yR9k
EyD7S2lIzJgW6U0LiX0dmYLAdAVzSOFZfbqex2lsCZjLxutbPMcV2d+tMpWFz85MH7BuF+DXR+6P
h0mohjPw6cOTjOjsPdtoI7I69zM9VWVHJKjQdkm/y07l4X/NF+s1nZWt2FPU9AA48mhx8+5KBNrU
sIyUkBfykkHtdvx8l2id/bZ+ixCclC52qXT7Fe9HMfo/1WS4WRq59G5Dwm1grVtPXgZ9tpZhY6es
kDCVyAFKRkoSDAWdjmvsU0lWcIId6oa19oaZYsvPYTsEucri512oB01CapWtCT4mIh1ND/dhkkfn
kq2pHhMjc+Ed4xnEMj1M88B2VmesaGTqpCuSReZVOqdt+b2bSoCHXciXR4z3dgz01L2Drg6xovHp
os523lSCpw8oJX6r/ElZQrDfdi+5zPXix3vog9UD+waoodgQINUxjczQ8hu8m24kiav9qEjlbT4C
Cfdz8yBjrjcZLmEjHJ1bUAcmSHhrHkO/V7XuzsCXyHML2H4J0X9RRznkxp/XEtnu24gJKedmitep
Q42n3Iim6Y2M10MEC2wj2C4CiAXiSxO5RqM/CSpv9e4ISX9HyPPwsiobTpLIwwlhIimSYhNZVGkt
3ABvhj2SbXIhDLu80XK8sXgBzY56CbmV8b/j4PBsx5NW+XAKak8XFkUUdeNpkRfel5vQtR0kSYiw
+wyy1W5z78vRKX1pMvBBbgwNq9qev6xWbnvPj8mBlj1rpg8IQCBmjzBPbG9o7MRn8QTl35o+LrxP
ti1yFJ/qJtsjoQ2Ona7O+Ea/+8x1BjXMWkaapfbUd1hZJOFq2rDWf5Zq1p5Qy2r1xGtPLP7Pu1Vv
uwcPhBLa4XWocu4h/kGkcignI8mT0ar7KITUphHOrrADusA4v2P6ajgtSZhFonPmsFu9dMRoILA0
ky4UdA3MJ+Mh5nM5Dhvj9iIQzQasdzipiSQzlQ/J+P89acWw3dDYufJUl1NlSnY61u13vaL+cPx+
U1wdHbyVZciELJNq92wISsje0VCO7RVBWF1bgbCuUnYT91G0jBmXaDk54Ibzr+KHBHgdXhTvVd8J
ehmq+28IWl5nEqOtaoAxyAvEZGutbzaUVYZyrQyhSd6LDCnzIJfxdMb7IB/fL3M0K8iHniIdm4+E
nugTqirnTA9LHyD5XNKtx3vq0hCBTMkmlTEUJQj0LUTlVjxdkJ0CZyvR/L9YbeKMawDRbg37h7kt
O9EvlsZjxlv0kKtgipNAW+JiFa8HfXlp2vXnL8bTO8ZeS5zXsFsFFaxbfzE/ejx/ejmYxborbNEi
0A8ldjJfTomUalpZ2Jv71ZPu9wpUJCDjjEn/87bgrmmm/i4+2h243cABmrxfb5P4rU64HmcwNzio
BuzePRkgraZ+z1z4G9bM9xP7/Lx5dRTey2akEajCZc5EFKnCUy99ly8G1746k30HSxBDvHAuN9VR
QHsO7+H7LkLVjJ2p/qyO0JZKqMOJ7AtQ+wfTxY/nKk6VizHqzBuw6P0NJP4tbPwjt28GMR4AWk9q
lZJeszHRgyOff7YyyXGsouQj9awM1GWiNbOxCxoYNa1M20BkvTasSjJWiq8+skWSGBkw9Z56a7iu
2DQ5o6NUxC7B/x+PXH/abZvQ4rhGP5qKYIycbF5JVoZVMUcUbRODUGPKnQYByiUFDPPPuUBNLFuT
aEugG6pd+PBqBjJw8ltWC/f3J+Y5OFith7dq49qsfkb3Tq6yymBFF2I4SCPbdX5RYhf8zv1y0dGk
oajYfL53mmn1MxnpVUbGFtQsE5Kh5amSwO+rLFPGLpl0+hPb16kPdG8ZMEeHlobrNXzeUMCVXCmJ
i9Km8RPTyE/V+cKXTehrORSCeb+bAI0CfQPl1csp3pmNgg/Yi/WGo8nElf0rdAQBlVvb6AvzFcuE
NRcDSCR6QwFxaxPcHGYev6CbyANYVsiRrJR0JscvI00zOn6TnyK5/To1GOgyuLUZwUk3jhoW8ov+
PlUoyhrjZzM0MHeAWsyjce/n31EQr6l47pK1+zWm3MmC6XpGLgHBjErDvsK3f7HMlqnOYLjvkPGf
HsvKqdVq8lE7VBaDXBVtkmhzXD0+8AEY1Tn7NxGGlTU132NLnccTNHRJkBx2WrguGZBYTvmi+KHN
pcukAc4LkVoNg/4ayum6nLFTtDUWL2dwIcjVnCvtqFVOyEQwWFl2eUJU/6/wHO9e/A1ckmfCbw5m
dEREd7d5LorEq0WGWbfd54DdBwkf5QiwLT8iR+fSS2EYGFIB0vAFie0NKLffNNZuzpMOZUThjT9P
SAM2q+689spERm9Ifnxw99nPgJFHN5gDjGjO0QJzD/OfNT6z+qgYoHjioz1ldOu63BsHhjUDcKwG
/eEeoOj5JsCnRD3gk+zbXgi2CeVJnJJMNRB3Vsw0Wvwxk2JtaU044ISJ1/ph0uYrose8iJGFDirW
wH5yaArimKvbVmESKxdavmz29h0TFKXwKD2hqeLzxxPdmFLF9wDPdtMMrkh46O2H4VLCdfIPFeAZ
O7wePOP+f+/toNC5h8QjSTfu6HTxJY3xwxXOO2qfPbULRsYlJ1381uYevdyeD5DYU16pdl6HNKDv
itbPJ6FYdu2ZzaHOX6Gs4Kw77ZTLbw79g37AaFpYGDQ1Kcil3Am5Pxl7QirlNhEOP3BCaPTi8mq7
q9ciPGWCEf3fvv/68qtnaBJXWSohCqC1X1OY0jswLjhW/IcmliVEx0qFbO5CsED8hicN2qLZwC0o
J1bTsMVUkKr/PZv2eL1FpWZqRa7xZPWuO4YfbsPDgrAyNewjQ1tScJx2njcdzRzQBbpho6b00GRy
LVDx3oSYBsT79BZ6rl2AjhI2Qu8MN2dma/c01jEaYxHhIUyKDzokRXUBjKIqp43UPdG199JyBlGR
O3acsPf7pffu82zCP8psh5Lt+weTMSW2rfvCsMcSFDRlAH7OEh8K6+rUlwbm/oNfbJdN3U14MvqU
zKhCxHgGM8FvvW65/gebUKOFDph7O1sG2gbE5U4vLuOE1wIr1krK7L1wSaicVZoFPuSFMtsdrdVP
q2dtqBfXtuG/cm5o/IrT5/db1cQGq6BD4bf5CLeOBhTeH/G/U7j18W27k8f6ItmMwPo8ABejLrZ0
0de81yCh9LtsAdQiqHH8BIO6ezbdjReJ2thPRWjldV/Jh7t7X57P1qD/MgpLSB043A4uqO5onwK7
hKOSLRxM5o1JW+Yd5tfZrVxbH6JSPQLzyaA+r3tOsg565JbT6TDQTuWfvH0pLVJjchcGNVHHnx/M
kZ++4SezSUf1bG0PowDQNW4gk8EaQx2rFhx/DpJDBL40paWgJOoZ9l0OdFBPD+yGohn1Uqje9gYh
BdYLbEwufsuFd1yYnlnAClidhktLteqcJOa09icDEyctMDGWTE469vfO21itLI1HiZMDoV4yiNWZ
ln/w8tNEYoRnxSGrrSiZpGne+9dqYPVfg5zY34gFNIGkl4L3luD7SrppCi756vqUNbzoCRR4qGOK
JssBmyKScSpXcbab58j7jgeFDZ30P8TZ5oM93P+S60eybyVG72xmPddOHfnKQamoYXAbNd+tdwwr
nlj/8nt2g0UQZqYtSyRDgthnkDMg+p74P2Yqo1tCuQalG7Mruvq5t1VZ5dMfP3ZLPPUBo230Y5TL
dg3pCjtk1GC64CnGAgNJDEa/uBpwgkq8q6JNEVpD+qsFXLXMayLVxt9g2ckSrGlvnvjKGVGpbFg+
TVhiWcrcfaqALCJ5zoJIX8nFlIK4v0d58P+tQDdUCLomvfN2ShZH5jlcHhXOWXCa6OeAvA/tl6BY
gSeHlEoWXN3OEH688Y1ycqYaigptXHaGutDMykRJQJmapdeHL1Q+sc3+ggl5e+LVFyLKHD8FJzEi
mEiQrZw/2un3s9uq2T5gUlsU1iWEDpPs4gOd7+nIL78M5K9ZLflCIcOBoMRnoYtEpceWpE1ucOLy
s3hlpFWJ/cUuStzUJuzFp+dAwgDPiiDuuln3imh1YrInhqFi+9Wm0mLDyjb/vMlqymkgKY5sAy+p
dYKCtmJaD2M83BjrnU74whO3HGlJEeoN0Oj4qjVf9hYQ6EsDqkrjsAm2d8SASlOm79fVqU/GS3SQ
/fiy7V+iOQfNhCXITmDHYKKW04pFS4C/wm6lYI03cSK2DcOXwInzFQwPAOwEZ33knYIweSfwXM6m
oJmpnTF1EzqLLRS8S1YTfjomFPtUaEizOTlGBPL+63ChhI6Obv4IuFoQOkKswrKBqWd5bMv7Ktey
L143A4aKsP6ZpVn8eIXCrzdKWDabA6rIOQjw161XSEVLyFjy40OTN3bv27hdbQ3pmjAdmajOrdTN
Kvb3uFBhVos0FJXNjI8nBAMC7fKkDGyglEwYXS5hCs7O1/5yNkNsl0cfaFM8CtOsC2CP72pfxuGE
+KMvvG2KbDCL8ZjkmDT5kADxrVJJeFYEfTKrHAOSyaCBinYzXeRMpj6+91YFocvnEN+p8CjKOHTQ
zW0vrRs2GxzVvWXNfjp4n/Zahv25BsAU0UJeR92ZK6dI/Qt7ZuZEpwt7wrzPGLcQSQrWXiBu0l5I
nIEvV0pLl2nuY+3i9UKSgnn5Aytv0+lUiKyyu+Y9tBD1Cbt2cShj7AGMExM9Q53fGpwL1dgVceLD
XWeIOUYyVcB4qFX22KjGefc0BtLgAawZ9ZngDlkGET+jg6WtKVDCXlo42GRDsfcs9/jN2Zuh+4cf
k6kaL+GtFlIeDDrffvPvq7BuATqrEB9m60dCI/f5sDrUvENMHway0OhfJVhJtf69GnWgY87VXcJT
GE4qvq9EEOivTpEsfZeKFWX8kuXHGXPQCiG/QGmeIrQT6tCAe+KtPVIXEFuUcCsr5yNxG9TZ7Atv
KJpkkxWrsA/TqDIGnefdpCi0a6PZlC9zT1bv1tduvGKSMdwS2Hg2GZDtJuve+ZV6viKFeyALgSk8
rOFpWkHOJ7o09Xslzijs/qUNHu+HH9hF+PfLQQ7kGQYUurnoV7K38Wz9IWdjrbdV43knU6LSwzU+
ty2JkaL4xeCvzyPUUWTt0THF1+flJ6x/naOtEl9ln8ggvjCa/Sy/lMZBcdYqmWniunwQeOiMrMWU
WppfwoceS+nh/kwyb3KWLTSqWMQPnBZFJ5AWSmqQiEVslbLAHTbdgkXa4qQieXrcJQtlqxlCIIGC
97xJnrSFrIJFi2Z8dswjsiF1fkxsovAu9Xpm1j8LxJPj49QrrHxSMrzZtwzeHYwBbduzzAyeDDe7
k5pcyDMxLIZpRW8NtihP+6eX3BTUyF6thMmQY/XQMstaNRAaT0wdSKF+fPMA8INaude/Qevw0cj8
a32NsThodEjfIHK3V0MvuGcr0rKR0KMv1tre5aGwW+FBJFwHYTfwVza5Bxojbs6iDrQqk7YtC+gh
o8Czkzr4i4TupElUYs8H2Oou2AQbI0Qc8gnS9USGCU/HNuBw37+MGqy35vZBb/MIDhvtHhBZEt5L
orT8P1jgRjt/66sVzzr+twzQj4aqxJ+NArG3DUISJbWTuC1LwgFI7MbKp6W5znxaadbkezkRf82R
nP7yRkF1c+zOcR/VWWn7pWl16gnLC7uyM5NAZfYoGkPy/LAjPAiSyn6BN+JwjBx8HnohjSDWkM9H
ddvYnsFzxJ7Lv0ajf6upPf8oFMxQZxvPUJp+t3dTYSCYZXtcm5t/Ahb/PFWulRKRMteQHPhi7Giq
8xVg4KWLVEq8bIzEklqFqFqT2eskH3FM2BIlNadTXC/yblCU52EbPy0lkP2DA+ECyDpr+FDlgg4j
e5oZ0ZRINB1stcUjDzW0OFt7nb/WENXQAB6WnNzgs3tTgEGTuIkNsY0YPrdIyVin93K7Qd7aX8nX
QLwnrtEM2AGl81Hltx6AYUeiMPycZPs0swM1duYJjyc4m2caf0+0VR6l/MslQ4OoWiStmYXLr5Ht
/M6VzwlktIo2tKPs2xj2j9iYShyx/IUqvkyZaJo+So7jTpt5wgYGv+2XOowzYTSKSyjIn8jqQRVo
y7ywkC0XJlPk3Zi4wqtvt0Or9tVJXxmBYG4SEurjSqIrf6wCzofqKeSEkQ8YWETfoKdgWi+G+FC1
07hU/5Vi4aKd+Jl/L4+OOdxqcJ+I9S33kwM6RUVakspk/6J6XEqLfefkcLNhm9f5ZFTSR7gQ6hBY
TvQUNzBzEIoSi7XnQyERcY6FzjpomvY/9D9WIC/+ZV4r4Tv7kTD5bCYJASCPUbOOvMdCHLJYSUgV
OQvtKzmYbfOYwBXz7UFd1wS5rlZjIIlq9PlM+xEiucOc/pUc4ZLuNNc00B4DUj2CqyQkEm1JjCYE
gnaHF0fXRHBBQMN+kTYi3d6YEYvTBWzZzR8BKHpl1GtYmGN8FPmkMXF1R/OtXSz3aGaIZpcPTq3s
Q8f9KRWU4e6ah6hhwzA0A9Yi/gQA8O53Y65B8cIKft1h2SfJEZz9wRhB0PpDxtHjG8yMZVV1Imj9
TZ9pwBqOewj3S0NikH2fpL20Qi7MdiWELmI/rbW3MXLXIHK70RqMKg3TJ/zobZrpWlpIRwiN4rgq
4xsUlsPVQRHgXwNVLx9jb8uCJiyQXDlvdUZw5IVgmLBNw26Pbbp0oroYqISaRuDEh9CG6hVPIR50
atocNv9zocCK77VR2kOGUE6d1w1xaUMXunJxlMM4wRsGEJGwm+27GSpmOvNFQPSB7NrpuGxRmy22
hIfNIIapa4H5o5P3bdNX9Fm1LO2xH6av6QACqsAIQqefQXTR2AXw9S4buB4tcT+WuCsHqhjxXK8L
JbdMTxKfV1VRnjOTLMv2MmsOkXOxRn6d50hSxXiUtPsSU+Kc0+7BQBhlk0mBLj/0MlQ/d6/VQ/W7
k9cNEGJVC25SbKjGeyOmhQd+cTC50jEuXMFuxA7R86zGD21toSi6sb3dRzSYVZcas/RhKNB/NYkn
yY3E34nFB+IifvCUxjXVrKOlbcfxa8pws85OdTmVPBrCIcpHYmxBoRVKRcJycWpUTLUMqj8f1cfC
1cRhwjKj9EoysbAaPfoFMKaHxgNVUvA2n4GsQR0MnS/O3NjT25Lo93GIsg9GcdJVIVF/0j9Iwsn3
F+n3/HK9/qvypGJBB+0Qhf2vxXpp5yToNPecCXTNvGmLdIW4R4lha+7CUzw51EtYz44I6gR7Qq+y
OHlDSUVjXNS6O3Lj3ey1XC2GGfq/P4m140VG8Z0Asik+Jmr2YInfE4ntGrCvjzRyS3WFIqW+UWst
ogf3RacGarrCiAQG7r0lKF3ouLDTYrrwrihRhletl7K2J/BXZq/IMPmOD/Cv/YS3WM3ahFeZG2bv
eetIGJc0WyAuYG3qDVi72++RBb372tx9QqGCfrX6hz33GfKsiEltAK7kIaM7VBaKpaAeyqHi3wkF
LqUkbI+7/PA+U3VgcdPcZ3CBb5ozS2d+11+aamA6DP48nXaDGtkHND3r//9BsjdimVT3KUo2IS7B
QVtOKBYav5UVTpTky423PFvlbwUx370Li7aA4HkxqnJj1BxwTuMuQDKxoovwZlBda7pI/mnzrUe1
g4rs/McM43qM4VXyrqfhBuYMAtv/LxTSA7kRG48kugucG8HzV80/HSxBujJ7tmJmotA1PwE5Et9S
t8Ps4zKrF+O1SrOHwliaOJQUTIodsuXd2ZlGlHJworocV1oytBwM0vdHJbiaZ22+jSppaLcC9Mur
NSotrMyK+GAacISExckhINCIBaerFEa3SGvlTNuioW2m6SBhSQC+vvBiu41GXLe3UIGL57FIcLgq
wK7nUhejpEdiAzcSM1gH1e9+HrozRqE64Bi+asJxNalxbg1B5hO1cMAx7GEKaSG9nke0srcdfsVg
ut4G5P4QI9GgKx+uK6G1xrkwayRgmqjYeVsRP/m1zTnsxh2IHWF26PpHVuykvvRZcS50qcIcQIqj
dMfXMFvLfvKjEfW4dsaYK/pJa82q3XYR3MrrMV2x85vWQcz7DedyP3GXbifW8GvYOmWQC9zNZAtx
VfdTC6KXzHpi9vG6j/ssmCR/lpraAy0OqomHhr+CUKYCns3De2UCmKZUlx53vjZxNFjsOwH/o/FB
KphQv4UEch3vW2EfqvEh4R8U2cUk1caZJCDM+wgv36Ix43g4xEsb1ineBtONJLOdGKzik7U6c2Uy
PkA0uPsKD8IuR6KL2omBcXnql4C2G2ml9o76sC3BAqDERbYDhBO/f0SXW75X+2Il4SmQe8bTItTF
K8wQHoVSJFfUv9N77FY8mWFTltkrFzW/6Nm8RVzkrgWOW7rJyO/lUdvg33ZAPv09UCEZmWCGhMRs
flIMlQMgP+YBdWBenxEpDYZOOZurZIRwFXM1LlYPyAa7ZzWYfPQH94iFpeAM/zI0+DO7mXlzbL3h
srurq74GaEgPI8zwCKROKCC4FMIoR1nwBwJvXppPUxPXejc0pyk0ROpCL7TfOzx9tIpLlyQiTRf7
5L1TlANgZKW2YTNGil9lKNLEbTcRc75JfoMWPL53W/gMYTZ+pRufZWmIc+DzR75ZmjIuARIQUWHZ
kdMivE41LhdE60gaERWC/6wIuH53hsKkO74ilgEbV+P1IENoubWTewtbJG+m5Z+uDYsIQ5YutV98
rrPW68K1uRSMGdoqYzsX69TYDmpV67ejF7fKToi8a5aNiL3F2+dxR3sBfKbUpc6NxnjYymbq+2pF
P+Jjz5YY6D25Ffna1Pu0zDZvr22e9tkrJin0tyfMgiPkJCGpLMzZVDHSbh7QfK/Wxkmr6AQOSze7
kazvV/Ju8Bf4THElEZZnafbMWTUXv5O160TaRlxCd3C5ZJfP5y6IeyksTjCXHoeD4anO6ZwUXPpm
941mAN1QaPvYwPH6N0873oqrEfCKQpfx5NDOY4UZLcUPq/CWOSbEi56Zjs1xcBODxbAAdOKcaDmG
qd+7c3UHO0i9C7ke6FPaDvD3AszXt4XARPvfhQPbvQ8RCxxJgHO6r9wWnMM0K1uZ8jGO1IUI7iPA
5U0ZDpK70RfA6YxYUXcWewLv7KjmJ1mJOPlTcoNbhMC1L57rB3l4J7VTQf33oxvoL/QJpuQFCjsc
2dLfW/+d/hOdrNf+L7QeiTT7iXkt+GTGFWjEnDAoVzNJ3C2Po1nUGkKvtdp00JOMVDoPKNMbbPZo
KRiuiZhwcrH1rwzTHEdBFVF6D+Ea+/XwYVgj4WRia1NlLuLSIJTlJSDSSFgOvvTUJaIetM6k+LAg
1EQIuGBG62QUwi8iFNkOUTUSHSJ6GLuDYyj5Lmkloo2tC6ytJCFNRLDZ7TVWfkP3aYjlzgsbRV6K
HwUsKvutHEpr3ugns5Fie5qq77Rv03GVAyA7ufX+a7dazjgXFvDuOp4zsdblvSaVaS9tgb6OQ6Aw
I7yMUqRYMqNS4DqmUteyXEf1c0WGX7dj4Ig18DwwsO1DVIRh2RatA4NxMjBlBdmOjE77iNG9fzuw
cUvurpqL3Mk4ry682+Fmo4YmbmQVZI4rU+TFsGvJq/J2E9BSgM/qyo/sIl3iBdJJMyK+/wFgojLo
NoYgpOdPWWVCFrn2qEAKsWmR2msE5cVz1x974RVXaizTcTeyppPWjJ2NXy5t+u3j392l+3egkBYk
eV4/3G51CxVP/OGe92ANsHqk6GmWkHMOaUsvJJhkI7QMTTKe3o0X3OhSVvdmyhiti+SvYubSDGdi
LUmG+Ni2zxN4dWnHydn3Uktl5kzEYzt6rLh5R4/1E1wbHwk/mQNVuUCUBVHLfLzzAr1b61tm/Pzz
Rbd/XZwh5kP0jiQC/YLv06hfmD99YDu9EvZE11IAl5WWUQIrnYQVRCxjwAnmOi6DPQsCdL/rQTxH
v+TRwuJI4tnYztIaZVsT+gynXu+Kcp6BgdPR3B4dMgBDmpHVAP7by3ntFu1cyZa95cDd2l/JIJOM
mrS5oJAaJlOvBjERi+dI2Ned4LPAgOtrUfKkKgNlROzoMpcogXFDuxpmcNHiAjOOmekCKs/YZEq7
GCmHH72i5AN+3X5A/VTeMYXTYT/jbq2EcdRX6yyJNmFGhCc2Q4hMI1KD3tzIhJfU/Ap+SoEGf0Tq
3EgaDXiH5lXNhssrwwy+ScqEvGKLfkMxL7gUxrUf9S3TKTgceCUM3AJM7F9grG8R5KyLHp+rCKMZ
b4Sqt+c8m8bhhziEAxBBe/5gSGffHR5hWy3zQ6l6zyqpki0T0LMxCStFzFd54I9DeIRV0QWc4y+K
mc6C8bsRaCgYNT6RF0VNff0uAx5QZcg4tE4dXuZLy/rjUCkgRNQ3WOhV7No/v8/9UbO4tiMYexSE
RjSTsDnlA+uevFxi4qxJq/r8ste9J1QTBc+OchDgO6tN57XkjT90vBCkfpaCUZp5PJKI/7qnb6e8
mttzh4vwCHk0iOJKJAVHmSDLYnBh4lCUFy39jbYsCEeJKhzvb3XqUJmVAxt9y3VdUBGByYDKEVLY
8azvHPL8k4uRYOVFoKjNlCYM3rXHUqbs1tX4Kqrm/1chJT5Q30faNMuyHw2voZV0w+OHTXtKSFes
bSaO8Gx3uXQfhCwcOcTVuKxhBE+aSQTaCX0ya5lHkRd0DFjhE5S43CH5flwFvbxs90YlbB5rxyd5
kqL7BNJh6vhEoPTSCMjdEcXD5OdQx4Rx36heNrBAgkv6izrfzxdcXB4J7RP9bFAdy84VlXhV9WxE
b38Zw8dJ1KBgx/183KwN6/Wa1ZLThl2eM/eYWGhu21m0l6uHt/whefeqO/shVrLY+YTGZFNBoFmw
15JgzbuAxxP83z1MW/Q2Q2/BMY3ELGOrastS9NAGcuI4yONdcIdXhSq2RWMFkekoSm2UYiMGUVhM
FflDrmIyHvABKRJdc22RFTUJoS7YmPL1rT4Z4qCNf5+brTKuTv4cmkWN09Hv400oBExhhWXWXfJo
tpk8R2RZmJ8rF8dxzhC4Sq4v8EYuqU25dcoWuoY6y4UK9HNAShuodGGBeIuKEIcd1nxL8izVHSH5
d0vAMVe1VANRRYWDT/grctcDWxMijCK4nxXYp4LckyuUKbXERWGLGZf619+lwLM9oXo1YZeazZqH
niaJIgH3f0oKHKzMH8mxbqhDzV3BqmUudPaqg+cx94aU3LJhK5hls9tWe8tRoA1OtSGl0bxGjzcX
7v3TbB1jooKKW3ypT3hVRgfJNsdzMU5TFsgfGbIVXKXUKa3eKK/uLVh2ZOcwo/huRGn4xQUGrwmC
TKaJ88FanMKUScEfJMKvKCwIkjvtQRGHgi1Y8j3Wlj0jPrFmdsVTTVdZtMCsLKfLtCgquOCq9bUC
uvEp1t90pkoS9PKnmPfLAtHkAhU36skPGSNOSCRSiQU5sg5mifxrA0N4vuOrw9/P07x9NqURRF1p
W/6kqdlitG7v3kPiLwkhhOjU3QZJqGBZP0+McBE6IWeDZ9ZGSMr+mbfZ9HYikRC/JTPXj1pm0xwx
6E2wH3584rd73DzMG+VCpRa3dOZuoVfmoRq+cJx8KT0t2U3BrnqMyO2ICt5JIdPSAwd+aQfiZDd2
OYTRTxPA8lWG+nY8vMBSztImlh4j6/yITyLV4szG1d/CapuHzFonuug8B4wJhdmIcMCxVcTlZITF
ntBNv+PX49k7XArYrYtFSRHssgoRHMv74EvrR7iDu/Bd4A/2WkDFZ7wPmQjR32skjdNO8u+ac+So
pW8vCwa/UWK91TNuir8N7+98cKl9CY39TzraoU//chFWk7xvpm3b1aKVyKvTT7bOhFLLluIqUXPk
qchUWu77lN57tSgHRBPs4Iw3KtTvClW0unXMue9JeTao2K1YsI0skY7Qit72DvytERK8oxB1j9YL
ouv/ndHnenyNUYxSau9nwpLbgovzKu65epoPc69AqpSvhO/slV87cTHkhX1MtOZcBEei8LlyR8sh
HlVF1A3nOLLKlny/UpwhlxPKEUpMXdCZEvVO2YAhVRHdqkJC5hiF1QlxzoOKBHdF1IYgXLvj3rSR
7NS6aqbOP6yqiJn5OQoBn2KqwrMlHT8O68RytOyyp7/tI8yeQgAGEjCT669GbG15UEmlKyOfLJGw
JYoesnpCowYr6tv+wMan+mHtU2qn5LHrIJX8FZg78MLKKOnj7fytkeI3O9LFjCTgYvGXOLS7Pl5D
bAna2qp/qecC+nOWrflZyG3wxWD3dEIJsGb0Px+I2Y2KotYhn+1cATJvCvQ9yDDcKEAe/kSMqlLC
cLDDoHJ5I45BM182L/0RPR5eDmMxZccWupo6LHKTnYs7JBOjL/g+N7MCiYiHHsarqphdOkSM95Av
Xga3lJ7O8nvhJ+btZUYiuBjPomQ/UlDPytPL1UBRNsiUMQFdOrWSxvO+y9jlQPnRdHso+ruuDFGI
/TiEMnas8JATcsfpDoAXqnAS+JJ0LeuwCRq4j12ZF3j9kLloBQHothENedNWKAbgyK4rBem6YoST
ukNSqt85T1Qj0GQ/9GaeQt83mIMAyAHxzXVsy01++2ShYnmUolM7En4zKK0BFsFVvgGdRiWZojz9
zTbM2o28fFdkt6hEA70YSUF1kKtNTvj+pqLCF1zAQqjYRRx9BdsOYp+MLHiFTmyiL0CtB5oV8uJN
Hn/kqKsHLAJAb+X+aQ1nx1XNI8Ei3CquTGpaq0fTQuIxlzjPh1e1/HfuTRyD2HlzkqnaFCH1ihfr
8ezKNrw3NmyIvQtQJi1eZtId+QBdkBAPFg4CpV5NRL4kZqvpEhA4s+vnTKuUYudQv/f0DNM5Yli4
3uh0OLH29bqXlOpHD3pC5NtJodi+MCx2awacdXkS91sx23n2kTXDnMM8VUUn9QEXm00B5/XG5B2p
fDjNf/dYqzfcDAWrYNy7ohPM3uyuStgUnpfA6Ry99OXvLSrl/L8VGCKDT0v5iz4Pep7/b+A0hWwy
rJ73MmaJwrveUb8EL6E5n86ZSXg+lTJCy0hgPXE8bqEE9wk/562paBh8aWpEjtRJUJFdeouS1jZT
KtMbfv8ilX06mZJQWcrl5cDiJN+yBtP9DjuvZfiLLUQ90BHhXNp9rrZmZWisX0H/07FyVviEmQ3p
DSxtuUjnWf1/ShcHvfSFN/gzAMNz7CDK611saTFAIEMiIbmKkpJbqMstjDTnx2pFaCaypAniC/zr
xMA/oIht75PdsORTlWk27I92qkmUd1a1EZ46OjR4pjczFHorYnbxRDJQuQid4Xc2IHLZp9RHQM24
xRToTdF+8uUNwYjmGVsFLzAkygYQHfWwo/6GvD4ThnCGQ6T/LGhlRMw/r4uzG7RNzGt7JOACus95
NPXeY6LVxnbUicfIMqRhhj7W9Ko5PBIDX4rOVJdHQR3ZPD7ZYI9AXseIOVZ8UBY2ruQGsXVHqujT
+ahVsJlI2dL1//fh+xQpG+EtlJ5OyVF14TyH/wJ2LG60o1vpBw26+/QBZgqWJpEkKLl12CYWZl7d
BjJzQvNb6w6pQiayvP0fR7G2EPO6FCHHus9UDPjXVObMJfOTL4OSwzxOyvbKqs1wK30UZO4yhF7S
zLqXjatihQ1tDrcmoypZSdr3fF+rdr7Wx7KyCaQ1NxwXxmY2DIHIWS1nnKugElyTqPxgRh8ECaq7
S3gJ8FCvsH1YkfcLp27xy02xMRlH4Nk6t/shL1QQ91S+jW+Ox4qqnKVPKNPMU5mtSC3Zq06FHp0o
yMVaFZx7/1sHoUm/If2+2yK9Dyt9HigUK4NOQgzzjBw3zzvdcZsF1/bfRNJce+3dNkdn8HrVYWgN
INaHF+6OwEi4USJCxBAZbRFyq/+dRbcvwN7fZWxJDQj32ylxZGSBW3SOIrVEo5OOquoSu4uVU6eV
yOfw5Q2GiVZyIR78gYHJa4yz0IaYkDIn01fGkazaalCNKViP/6fpOC48IiKgBDKLwC1a+BGKSTB5
saenLNPSk1jx7KpJlxxxNtD4hHjQV1l/aGK88E9JB/QheG0oLyX0Efx46Xzrpj0i44omJLXboxtr
aSQVosITsTd1mwlIAoatEZfMUK8+TlGbfKjsKsCslsFJ7dHn2sOZPTrNrSc3/1OYx8I8M/SDQmU/
0+8QPvXZ/rXJNIpr4HdQzVS7YXx9Vn+E+ko7ceVE0KYem8hIM7rTcip7x0TJA+aK5fAAZ2gmimlv
nFgGs/ETWvIorpn3jcouRRSphuAPDnp/keeikkjnvIzMB9MBttfn9MfPL219B+puuvv0j0mmZRT0
00f+VdR/v0V7nRE7t+y1s/oWei6mt2UdxHuCOGCWMzLMargz2cuXhwxyFKSjSONE8D0LGOidE54S
JvvOm9r0kGxMllyWXc0LSDDIxhIPEJ9NjKnTWmf7YrZWRoeKSKyrkHZjV37iTF6RB43vQj7a4IZD
4xO2mrhyhFoCZmUsZD3GXbSIn9UsIlHeXSQASfJnjlfFDCOtfRs1IVef8NbheZpBl954xsa9bO47
qvopBo8Xq+gMG7ZG5OYM2qBRIOJfPIk3p5GWP3cVF6Jb4Hymai8qC/W9nZYHvAeDnXtBeNXfJkA4
LmbIg9YY47c54O8wh/MyEj46dlQarPhZEM2a8OZMlUoGzR2XrpJvh9yE6JspMfx1wrZlNCrrwB4x
qaykOd4gNoJnKvTcPtHk1ht+7+ckT9Hkp/qoh3UdZCak8HO1NNu1jb+JTvQAoCBvvLuIQXeBvYop
YTgAAA8E1IyQqK2pS9U8TIe7PYtX7QtQNNpDDp/8PFOyZ1x4dKbuI0CunUXBq4g5m3iahXggi+dx
FmypL+kVqMHfFM4MEmrF5v4kbQLWSaiZrLW7rMq1nd15NuYG0NIvzVG3j3cesMt1fgHwK3lJ81rh
5dCZSpBBLu/h/KQBmBiGrcb0zlwQfDrq6JFLsJn1JlkeajCU8oiHygEkiTfvcP29y7o+0r1Igny4
si0KmoNNz9MIxbkRmPGuKeuyAgdu+X4Sq/MKmfRFXX115Qbri7pnMGgOSdAkaYnMe13W+rBX4agP
kYy79FC5P92izo4wari1vpC9ETSVOnw3IAUYyDYEx7PV/KIiH8GbJqfL1ypMCrKl76l1lh5pVtBa
MeOBwsBFSlg//rzXX7MDcxrb5TNDqk7JehUr7a9E6qdqSghCO5O+GE7xwawK9SdJqdjX/2rWFtEx
3PEPEoTO+2LhLsnuz4IxKaK5ie35NIYRquYCJdFnQkvloaRjzL5uDanPLVPk3kGGWnfAP7Y026XI
9JcVsvJza93iieGhfaVGndfwm0+/13oUv0k4V84KoP1nSdtZ9X9W4nZnxoJVBowPoAyNH5EtbzYI
L35LaXfyhQ34Hr/DCyGLrdnx1FCA8MvbZCol1HIyfxno8GqhUaXYXWFaa+ap4wprEJMz51dz67m/
3iE24Kpq7ZbWs+Gf3UMgrz9Fpc5OLWCG/5/HalQ15G0yJoZqISdd+uzvef6FKr0/zTl9s0lf76/I
cBdXxSnymfc1WmMETidy7Ry91IBZC+6ShndGC1VYo8R2QUHWv+UN8zir34AeYCB9d8ouUqZx9A87
P27XZO2tzZXED2oFq4b3KGfTOa8xeD8rUqZTM8T2Cyw1qwcFQ0g+PncZtrPgmtr7iOF5cAcmYfH/
QOZy8G3Dr+MzCPI4oIL4SDYR7x2vKbD/rIAZAiSYwNUcmeC56K5SWRnUOFlC2v8/l4Y0Si7CS2nA
bEJ77USaBJEO4GoozL56sD8GGkxQ1nbdtprQsOBLMLgVFI2IaDSs19DlJgnWwi31XFYrBiLd4c3a
5eZdj02PCXJEfzUj5FJlIIy82jTMRVuEv7ZUxrUEjq4LZ8Y51ArSE2efUTbHOA3frE2ay7/NFHRO
b3nx4hQh9t/DfcyYzIV3nQoEhtdSY1esYa7Nix88UIsUV0gZya7s9L5m/5JFT2MTQgIM7caaug0M
vMDTCG0zUz7/kfK3XpHrIlfh+2bs5/HIhbx8NwNwRjCJ7lewlcW4T26odUTJwPFl47iLSjVll/2I
VPKXdk1xANVPK4Ls6+n9J5V1P+nnKDF+6NT3RI1kNQx6TW+tY37WMKrqGvNIy5T3vcfHnHKinl/S
EfE6toVpKfgQqbkhcXx4cGt2ZdeFpiGe9l1J4xywMysXh3OZAA4sQoIW17zw9HbmGla4pZVDtNBw
PUHvKKYAcJcuPonXduLr2bA7qvHiwR/T7/+K4seusBUhTrbUxhXwziSFNT9PZ77Bu5NBkSBMGbfo
zWXhSd22XpCv7IS5vJhGuMGGpxWPLi2deJj3zxQG4rv64wm+eC6vXg7PlHPQ8KDmW9W2dB8zq5yD
O6y8svc+pOc3bLH8Vw7DFJUsF7SmomLWMupX1DUBeNWhU5BUYQ10INAL17A6isaOCSUQ+kgh5pxF
PmbGxKzN84VP0yg6go6OXh7L5rG7mBDupRNcx5SB7KiKt0rKRr+z3TGuTnGLECYd3h1fIdA8vJOV
t9/dk3qxv0BYFYK+uxhnLMOg4q2jbgLZx6srIBXTF7fnyC0c0wFpOXk7At4K4th/kIRggBIy/LY5
i9Rwl8y5KkQubt7ZNY5RScR7iTzSMbnHCIiNDlVCdt6RvHE8pdnSXi8dzB7v8tWVOFD+xgcfgRJJ
5odyShF1rZVoqHEF4V4HD2Qw30VBIVFafkZd94IILGELN/lpKyMA81ihPbCXUqG6qy2DTnYmTWSE
nCbLTkQWPpCxPM+RCSOSECkZsjak2VCkfSawocc5//xydgVQc3U9r4AsIwEaMIZtWwc47ptAiREi
Fo8HKolXW/Nxgix8O5AITIGJ/J76h2zBPhChkp8pD1d8yWE0O+tSRCdx9P/QpuazyfFuKaEH2YXW
B+1bwu7kp/tj9xgx9mtvq8Dmny1aPywYEidewwSBMgKWjJwsKQt89d3J4KuAtP4oeMoeeOf/horJ
o3rrCgbiKHJySwdrHYs26HAR8Zza1KPl6crSahSBH2tsmXxgqfnHUsGLUtp4ZMA3BJqu8v35O2Oz
AmGPR6lUd7sOz3d38bTUV8eRwyf1vt2ZWajX+qqJz9jutt/mjf50NR/Krl3M6EiEzZPKR6qEKLML
D5YFlgVnV/RU4jAxxlYGp9811uqjsOdNe44gfc2BS1IdgCPKXS4Y6ce9bsoB3xUGlcu7hDxkGtzP
7x/csCVZOvBOMFfgoZGpxQrJyJEq9uuXIp4bKo/laEECKEfsL/Nazl/F2woODdoECrkjDeBESYeD
LYaHz9wUSzr5yIBnbsXXY0vUYVnEThzPL4J86F9Qp703caF3MWj2zG0fOqwLABiTA2vvPh3/hjUd
7HN0HE7TzbyS++mnW3fopdRFySiMS9EPMoR0I2H+E+MkLBm+HhymM2kRkXwDdWiOkDFXnHrEbKjZ
vuyEu67YP9pX/h1ftSh4iXE56FEGxi0LMzAnszZ1VMjK9uOwe5mS07msHjOMOJXH4B4TbkP3Akkd
KAirpb72Db1eBux7r28u6hCEsZKdgMVAS+IcQdTVoDT9qXfudtGszK8nwopN1Zr0YtSlOCIA+iS9
G+qCIJA7eU/K2CZ/2/xO1ZBIG7L3gb7cJvI5m2p3O+Fmgyatw49vrUjs7AzCfyAI8PXvO7GCXGKj
kh89+3tE6vhku89azFpshr3sNnVFPulm6gshEPmzhlg2RQJFwzzwl7xzjbVY9C4HTmrUZxOIT29K
uJwnM2D1RfMs7O2vPwd7Hohg2VYsYFWQoMqsRmFwyKQHQAM/ehcQcjPn+qSCAoxLcce9t+CZHOiH
KkFoQ8tJvtK/wlTW0AyG8dgy8ZzcHIdwoOIprl7FMMjJkzEO1CKLA7oaqU40k9lM9yNFBDlRQfaV
Nn/uTDJbGAoM+FTIvDRXMLd9jcsInAuwgxbZ8lN3MmMlWKRDwLEszNJUTBbndqyCnPWL/977sv4B
Uhj05YjN4jHCse26Y2zz36MtvYO7kYeqUV3yYFTSN/ZeiWAi6hUmBrRAGG2jLY8fO4tJcGJVDKWZ
ejBkKWPY9DQuFtgmvesS5ZNtdPBZyXxUXLw92Xnenl9b6deW5uK1LkoDmypM4otOwIZxUNNurVeF
LCjbq39ROu52r3gicCQaz7g1UcNc9RQgDzGC9bi+KlAdwom7b26gSv6glSCfrj3jqSEUT8Om0mfW
DyquXufPnS5W2Rk9SnfuhZTin3SIdT7sR22atimozH81GHCApPvzET20P1kivqokEEeFmzPhC6OB
KBUCXm7Qjd+/tZLiXRTxFKI5pWcbB+YjMWYNGlu7NTfYpO9h6nLoP+gsdRaXuUnY+JbUhq0TlRjb
waquYuWfqUvPQ/Q2vwhY7dHi6p4sbYR2wPVAIevsVDa9MGA9Zhxdb0/BMlPgUlUgX7TIR2vS7zgk
pG4SlfMvlPThyQDNY1PJY4Rde4X+zVOO8jP/KzZXtetUjXpHhUWytluC4ZNktnD8rIwBuVTkiP8w
9TvDA7yBUCGYUVZOpUCUubmnbPnZdBZg7mV/OMm/x7nGRXNmpg8Zhk5ycijdNRGTO3OqVaOUgbBf
vkzd7v3t3d+z5deDpN239xWBHS0mjn/nghhbDAe+NFuyFtuKJsFANMAh83k9Pm18sR2nMxrsiMEo
yjYgRVNWAwcewCiGEOopYbwh9n5DoR+CzN+bdOnMUBbvmbppNLf1/4Wt3LW6VP+w5D1qs4Pr5eQH
Elgd7sJfywZTmjIuOGuLSS8qSMNeAoJTt7E2KO4/hPUScYQIBZFkHM8W/MNIag+e7Qa5Mkhc4qtO
NWnqW1cwEqAD4sYwDGNjAwOMse8nI5P1u9Tp4w1rAZ/cFQXkZzFJkJaiW5yhmH627neK0oImA+jw
/xMJ2aO5bCWqYO24lZLhW079zhbMjtQtNTRwv1r9CGHHLN8KogMJghbx4yfxckMUkhPuYNkh9fZP
oCs3EioDIuKoFenO1UmMegI6Ha/rvYUEGZkcfY4CMKatDa72o9QxWqvmNUE36U9j1cy/m8BUsEey
rcwvOykSjHhI6UR+aIzeEmEbQwRsnZmys/E51OtpLPo02sFB8Z8QXNwEVyQ+iwZaPcmr0S0abbLR
5VphMdHwKs4Ql97EoYFArb9AQpFktPDSSarXnr7XIUzdSs5Xq9PImUyEMn4PHsk/tyIdowwTFilY
gLKcZj7qFheasv2G2bGlKo+bdNS+FmZw/GrmN+Thzk/EnJckiaUXJH45wN6Z8wI6PtvDkEinLISu
R5tpSPvCbv3pEBXygJ+NmCCU7tsQNryPQw7d52AsVECWXaYJBsFhQc99NSJ19x306EM5SoW0jX07
5eY0DqbbYfpa5wZS6yxLc6OdgVezWzqzfSTi/EJHUO4VhCx3JoGuvrCbHIZR4cJfKle4HqIZeCt5
FC8u5kFH+yRv2GvyCekTM0H8T7q1IBNsrbKvKrjjk9MvFuDHD8zXzpiEOt8HFK+MnlQ55zF6oUBH
ZqJmJ4JOaFIeqO04AM4wsNnX9UbBq579c3InNiy80pt9i04uTXa6Q0OHWZPbPAYVimR60oLw1C1Z
Ld0Mr+4fdYtvq8zOdmiZ4BrYJcvUbZ/hPG/yBSecCPWny1Kk2spYD/mINosZNB6GQpKEDz4QsO15
K5ztu40kdIpGIltdzYHdLRIcTc0yd+rSb7HDurYTuMknQ9aTqaM5Ee7OYtzUqjwypE6qxLF0C9sZ
9Rp8sOxFzzPvKOh4s0IUjRDFXfEdMphOlOkrUlolHfJexzaez55/vUI/CmnUlhcRENbE/HSofGAv
YRkckkTwCLhIkUfty+BhXawYyziC4jzUZH9lK9Q4hg8FFo3GGIeZ3Crg5tfuC/gSmCtrRcmAjAzi
6RwVGohP0hUQmMpJu1Qh5qrdlVTn3bjFw2o8yiCN06b6PaST5QJ4tMvZJP6+D0VWdU5n+UDtxPze
FsnDPabRZzkimb21G/x5rt2W5MuMuOigsl2Hz5R+8KyEfsgn21IahITmJLfqKqohh/ijrLQPb0H6
5plqCO0j5HcNqzQeA4MnKl0t/vVrayXAp4oByCrxtwDpIIku5tWz7pZbw72W+lrH/pVvbffU1mMD
+Zy/l/ZruyTVVd7NkYYc01Pq7gN/nB2aexlNZjT8FTYgA2OfLDET7WDsWBDAPuc9cGbimKMLVZwa
5kBgx+iIrFiaftjPZDGNk1LurWSeCy9JW0AXXFnElsyYWb20EvHRlJlc8bD4hxJ8ssN94DlKbmc7
vPaWjS138okdkqGoY4S0NpSJdZZo8tMzmK+PTHzwa6jS/x21tcVgV8Ypa2ESslpQkMWJl+XjKFM6
puxUnH/QrR02xnS/TdQNgcV/jbCcUkZxcPxcTUU+IRDnXves61nFbZzkxDRvlQUtXLCY2UZdH4/P
+TjCzAnbD0AgvgCRsRhF5bEXQqj/b9/4BblpBCX9STHixmIoRu2BUW/EAo11kvTZl/blbFVpLD6h
3zutyLK5ZKWOOIfexufzHCrkXZTztVuRfUAJ2ai1CADB/o6XGU9QpiGoythchwpQnSjte+BlQx7x
fH46HRau/1xAiRx3q2gve1IYpbeA17ewXCYsC0ke7hVZ6emMXmBdjfEGaGQx/1xIwfpvWHwO6TkI
6gKrwdckolfe+trKy88U5iQ/HoCLKHguOLRZyk02JQAdPGdjqRGHraCUL60Je+KmiSA7k/OecWIA
t9SWKrHIFse54fxMlpxcbXFNX00wLkAEE8ooYpqK+l9HPFCd6kuTfw732b1HnqJFOFTQvHWOyvFf
MDlYZnSnIE0wiJjFU4ni63XE7Jsu/1PkWW0kiBf8vgcTeXD+rUYxVyvDgs8jd1WiwqEQfyKGqJ1M
t8ErSyfY1sBBbOdheaX7s8/bL7innkTxjooI26qCTX8RHb5q8rDSqpaexBacMUcudAfdlylweLqK
btc63ZfAcloby+KtkGviC9nxVO+eZXfCEDFBEYTwhOnOuTdViTiqMnjheyYoqPG7hc+6jb4gXVyq
pdmiwOTjCuzfrAhjolVZ2Jcxm2GnMEYnlfS7Tmi/8xmcnkeHS401qhhEPKvEUrdOozT3+PPoxy84
9Ranuzb0OOukpNuN7iATcxluM50anbz1CyoceTI1HZqDv1F8eq+SAZhByxdiezKO6kFTT+xwdR2c
1V5yq0JO4lKhFjzLRzaueHPcPRhKUXotJ1sdXiNhaAvFG5YmUlOOz/GNttQz0qLfPMhGONk3bBh+
fD88xA3dqVDXunpmG1XVTx6xL/9VW0ifUGqkfCpHi09Pc8NWmEuRza4EO4Jws4OgTj/66fioSv6u
uGbd+o1HXMm4opmOwIJbFX6X71loWukopNVs6o5DA0YBoLPmGuYi31WUI78r4dhiAFzpZmRA5p1K
poUtNq+D6xBqXXX+sZLcF4wvn3G8CKwuBkhIG6+lBwOtvPoPO6ytcD44QYL0yQBUp4zHwduVILVV
zrXcTQPtIeVoj1D/w7UtIgyQsYM3kx5pA1dFRvSG9ho+eyhhhy0044BDrJO+I8/EcyblZ2xUwaKV
tnlRUuWxhzSQ/K+UKGVoSH1fL3yiHGICgUSis/Vd////yFhM3GnFS87xprpetfMYmxeYm7BQipC/
v0vw8wV89bOjjCqPfG/Uoc86zey1p6xC8efCpECAT0lbip9p1F/4gYFZwT5Ir57jpvmheUcyxlfp
VcEEfXPKE9G3bpgxHCI0nqQj4OAG6Zrl96UzCTQz+DR9vygDaFEuJ4M6UdP9SFLtaDnsQFl+VMJp
Ej/O8Wb0ddr1APh9z/SH64TlTs9Eyld2M1o60RpusfY8sz8OBo9OLPH0fuk6l8bP8pEQiO7kfx7J
opiQIWSgXl1JrvATsCanqUX28fSKyQw6qslfNQHAOpaW9ihEPpTk+4RnXNY1XtFiSlC3ZwjZKP85
k0akxE2umlKDRg/Lh/3OLD65vvj5k6x5zw+RuBi4DaQdE90tpNRBGopxa0pXusLGljECQsnadxbM
/c2Ro2PrLDCuEp7DfWhBwLHR4sv9qRUBgX/lwxAeP9bJ8fMiCpGH3cQQOsoMFdi9hMZ0o8W/n9Y6
bpDLKPPrj8nIsWAJgt/bOdhvDaDZm6i5j7HGVIRYZ+vNSDdHTL5RqSxm3vTw68Nd/C0yA4tb6DNG
lo70WKw1jJ1jTw4eHnmQ5J+pdM/iTgJGFJgtOJPDumeh52AxGVnEIxRUR2U/pe3k5S8ONf91FlNy
jr7ya5KTQAjaDKoe1WkrahTnCcFrXQa/uIJCDAtVH4sE/6fa0N9G2q4ZU771ySvQwo2UoxLBBsfL
ej1FoS/s9Xwru+APZi5Pwg9mWCFiOa3BBTsUjmrAmYxZBq/2bx1M4LMMXSI1Br+oX3f3CbQErQ23
vmw/AIUnfB0LyKu68UoMDH3HXYE4LtUxIgTUd0svP9KoJrlQvAqBI+t9oNsNoSqge40jdSN7orr1
E6Fnx0vXnbcYIuC8R8M00AyreaU7ysIkgdikJ2gYJZb03y0kwN+N7S5s12duo4sv/r8qeU9aq+zm
r/k7f0ofisxOCXlr2qgwQLgkAfUpIh7m0buj3DTSzdBrEJtVQ9k0wYM+Xm6eCyZ2/X6W3hXAmxFc
pSXeolq4VkxgG+jlVPUMSGjBykcMA3isOP4pIyvvPdWxXbwF98o3o1ZfifbHzQ8G8+U+4lOjjhBG
JNLT0AfejTGgmvddF/8UlaoONFcdt5R9ENXYZH9J43Ak1fe6hWFk6qTrS3HaCQw5uenQcKj/Dd3K
U8O2b+TtJrIxd4PMehbMiLO/I/vgYUqZcaBi/cG8+l6eE/e+1FSF1I1ZCIPP/0MJVeJr6Ke2bnCQ
N4KeN+nsy0kwWITJisgDpV/KLoC7GpYtVHuiIrEs9aIV12ZRlcn0TQ3nKf3mU1F8Rm9HxMcmfJUX
NLBIcaqsvcymXj2uP0Q8b1qBWcpXS5nyetXkXxgFAJIzMspEvQLcptlVZpKZ/whDp0VNlJA8wlkA
e+bnrt8JcD+fdjjGVd9QYLPat6ouw8ReY5KNlljNTP4Ijn2LIemm18+r62mhmVxYcP/JCWvAgXDb
rIA0UWtkxdos4AlaIW0Ts7g+PVopji6UnYHWGU8X8bUwgCdv45kfe6hCTH4CVi+S/MaukwlrNaaF
MMLSgim/Qtgt9pn/rDaVn4Rx8kxXeoam1tYKQhzHG8Los5YZx62x1MGGXT80eR7ix+3XEOcQZmyS
xllzk6YpZgXXzQ13ikpGb9Yjsm85Sd1rUsZmSav1/XsRihUb0tnNG2p+KCXiUYiQAxK4+TobS5pM
H3F+lxqXGdZEpatuK2ZHtliInb5nnW5/htvtDWikclVepUvnR/JBfEA1WF5Jb8F8A43zIg+mztQv
1N/t2Wg3eXpyMBLKAJPujjw22ZGwEPUTZDIv844hbX1TRUyEzDjFO8LzEvM1I43HIACO1hUK4/Ms
ATaA9LfJiSxL8V1WyuKOMEULDGZiK84TLmTV7zJpx2QZcvNJ3SaRMUYdprf1mNt+RlQiylJNBOGI
Tq330fenZchvNHNpOfwZztF1+NkgW6pAFJcBPnLkWZnCwq15+Zj8VRAvS/qKsyBLLcMyWW64gI7R
x+H/+ZbM1N4nMJBVs702yBgGHXd4HhC4JuYMJnYk5nm/CYs+uwvc8uW2+6IicBZ4Spg++hkOHQfz
ygTKUC4Kz+FU6VSknhUmkA5FeCgmrPonZw2Bq8/aWsf5BMWw/7XSwQcZhn6sj8FBo3aejyxP5yNJ
5K03+E5hZUDqGN4QfkBbA+MtC2vsdJbLo3CTy4g0EWupVIoFmEvndvVq9m6fwBlTV67GNb9uTJh4
3MNfwsnhrBTgmYna/h+is0DmxkvKoh6ObkVVzEOulJVzfDq2hnUoHiMI2qyy6AmguCXhz4ibuvrT
Sb1LH6r0RICOUxQZG+CNUSNzdcJb2Cac5uXQQTfsdz6NFl2PcP3l9ffKQylCvupUgV7Qe48eZhIF
obde1LtAqCVaoiGBugQ94Cf1ZJF2plQYntiZmr9IOAgFV95xc4l2sCcIlqmQ2k73DlqyH709Qmwa
sVcF0rSXNBOw1gwvYOzlVWd75BbyfCalCIjuFL6WaFfV5DXFP6Fwuiz/fhvcBy4Ex+4vUedWV5Gx
UP/WL+/CjG7szZ7j42qPYKZ9aS+b68nx+LGVDjoBOOi/j05YvkkB7vvXkRZaTAuWbLQJlmIy7wv9
hCTJ35NMme1weQ1Ga3PsqnXFEa6Wr40ROmG/Yp6UQAx5ZdoHyDKQgj7BjKAQ+gOATNVw/2EsI6xa
tYA5LUKLEd0my+67WkpRhpN48KXnUVbrs7i9xE+oy5FrJO0+9eNG1I2PmL5uklJTmPEGJhP9jGu7
Z/3pJunru5VKFTcJorBUfpJcZ80Qqgn5YLMhHjk3CiiuH/MOi3aXdeb+HQo1hMDOsfA42DYT3z22
uXB1/w0pBNmVe5D/tEYssIZa7Mr5XK8HhA12GswWgEMrX/BZpOkbZkn7weMfHHW5zI4eCHuS+6XC
VMHhIajtdUmgCZA6xcRxKsUCxxO+zrTDkAlPX240MQ34jLpz9LeaBrFf953K7/WOSRU8UW3WGGG6
EUsD7xKx3zJ4YaObKDEg13v6fAhDcUGp/2I2+LGiIrIeKwCej5kzOsMTYAx5nF93AjvTGu4AkU0G
qAyVUg53yjxIlNHSGw+NgBo9ccVWln+BN1WaxA5FC3eU7iyQv6aihsxQSTzKsdRlcEJP7wSAYZ3J
liHoE6cN/UOZ+SivdoTgj/3zCgHSK7XBAR65dePlDPKWJFPZSik1IEpUlhJpMfYf2g+XVnhXc+wK
xXPrOvMpPYqYPprQgX3RMk98VEtzaNbLKKSps/UL9VxT3BuvNEllUjN0/VFqxAjxrPT67DqesW51
KpJtktY2MzIDNA9J8yJk3KDBItHnWpSdsOHt2yw8FcHS3eNjajwMzYUAg0AvrIGqjnY59nMkfNlG
1euN4fKhkc6tofWfQCNbFZbgj5M7G5VKOttMg3UYJNMJJbb0WgG2UBozYMjivP9s+Ek5ddPFH1B5
vk4CVOvdKsmiblUWc2CE7jF3H3pvpRjU/C3paUz0jBbhToOJ4m0f+G4zEDUpDjkvyS51egtTTc9Q
b8/JB5OEBcvwGnw7RjpeI0gPRtqEpdXraDBN4QaMFW139emkUla9zVW6KscdMljH99bbSYnggI6+
fRxvPXvRVqhBszRpv/glAb0oTMdUZ83NiB3uVi6nk9fligD1PLz3qbu2/gy2TSs46j5UObKCFhU5
CcaIARzSM2xEz9ZTRkSSlidOSBAjx4hqdsdXDi/nrVT8nQ4143BBhs807vZQ8D0VvunE5OziIcDS
HVVYjeLS0MXAQqoaYfEH7iXvDWQDDAJuYzvBf3LwsY3gcT8OOG84BMcT3RHXfxLmnDCTXV+PRKR+
8yYhF7VGHz4tpeGKyUcGwl9Cp8YwJdaMOJLkhLwZLA8aK4/YA9QMc9LNlI7izPpooJ32xiAvX26a
I5GPJvFYHXo90Qd23vuquZlDBJCkyGZYLTvP+5KROuAYYKM2gdCEkXZVw8/OLUb6XVwjkyxkKNif
7sURaAR1YgraDJSJijP5X8vTmML+IMLPSBET5kK8+Iqw1yaBm89fhOy8h7YQUAdxDt73OzRBci3D
bJiHD5ws2pA6Vwldcv7bY6cU6DKjBpmRuOSzPbzXyOjts+1W8QmG9lOFNQAFa5B4Hs6+Vbe9k/NN
O6A3ayyBzFZ765htGzz4tiYLgkMv0rDnPtxAo6KkB825Pwozsd9ltwxicP6fzWube9iy8JxpgyMl
YcjSBfAIVrWGeQ+XE5JG1/CAL5QJ9nC20WaAkkEeg++dFmCCNUUkxiwAqJCwT6ktiuPry0wgdMel
peDJAQCi/OB/nEY4lubHYwuxDpz5ISuu+o5JO2XtRdSeboPksJxYVcarWZKkQLk5OgX1j4m96W0A
AusTlUfdGYRmm25p6lFCknrcjrq5Rv5ZViwo0xaUR3hQ1PsFeiiruBKfyPs20lGn4gdfDs7ujRGi
x72jJShQNkkot5JBAxPAb5nOaCN0sSgLG4i51k/e4TTc/8gjUBjafVlyoNfGFpfNwU/yB2a6mPxz
hg3hd7H5ROwLgET+nVxly26VRzMXtmKJPlVFIrQtaeNd5eHTdATpvdZ5/VX0sO9rnimKdMPn6hwI
sCgAsOaGNF8zGjEzRZ/2uOHnPEDC4lbWCjT02nCbhFES78Tv/oy0CagKO7/1WkDknZQLYebTYCQ8
N3zvKHlh7jiMuEN8F4HBNIChcoJbEByaUgMd1baerY3LLAZ6B1GjCgrwvo9o/OuHEHfYssA2vR4U
RXcIjlxEHnd9798s/wNLmPZ2vhwKb7p7rA14dYHA7VAqDYQ0gR/nI5yfaAEA6epad2xA0Ix84PEb
JFrALJg9obKO0hbqLpe2QXrJIC5chA+x7AjvDfwOEvX6f2aqbELnSkBGkQi44rJGuoWeAFkh1Lz9
I2P1NYL00tvJdDOc9KMeVeIjr3OaHGzj7qVWusGxaWjljbp3Itudt7Ej7opWyjVkfFMGH7Vnd6L3
BVhkmxmZ6U/SwVai/HvBzJgYDxEeSK2J3l8ofvbeGPRhNImzt9UNROoykRLQcWtg9/TINkT1at9b
8Awr7FyUqIK8rh/hlZmmwsmudijDpsXGMOQ3qFNqMYI6q8HM0KkwW9Zk4qhiYUYCvVea1zPGweiY
7wAfcPCay0Su287+MpvUsCjS7o0InWr4oO7DYAguyp5ZuChWwTD9oWmem/XpFfqIlL23t5p6TlOd
TRKDL6hReemCPq00QinAANJvfZICZ9bOFDXK/M8bn7giYUWnVEZ6ksMAeRQZSgXe/HpSsJX7RHfR
UbRi0aA1Zx09fDzOSCaqdvJItMlifOHqoLBQ31/dJOUDrN1mUC/go6YEZAaKc/5yuCUwWUPrfCwW
2lKRKdLCrDqDZzeV27ebpg/+dGSAVvU6Hqta6HNWoHhsWBG/uGsGTL4iM6Y5cWEVL3xrTXOiRU4f
1Zy65IqxEOHwbF5/UtfVbsspM6JU9PCuQzGzylqRvYTR1Lm9+cjsC8lx1PhIvMHBMi7PJHxRyxxM
1cNKY4j1ajscWZCOAzRHSWUvupDBa9JS0dOvjaB6xpF4GuH06k0IbTIBaWr+FaYzOnvIZCEU9A2m
gbtSN4lN7yX/HBetsZ9Mo/WQQpOSikTf7iIVf21yLDEfhJ6ECIdNeoTwzFf7aBahFpphxuqaji9U
q5qhtQi9XxQPMiiUX24jNQ/bv7ONHXVeAJn7wR3hZwhi2ri7rSCpyMkRe4yFZUt3GNADGy7YFbIV
tdUaf4E6zrDDomJgip3lY29ohgu6aY0XoQaPoFkeuMFsVUlt62CM+evVD6Fe4ljfYRG+X76wrIbJ
/e5U87uZOiSMdCoe28UVUHtMGWLCB+lsx/Lj4nnbbX0UNSZXl2U6o9MLaDHHU3dymGuCatmbeo22
cxwXvJ+QO30/bGlaWKQKA6P3xKRn+gApVGeJQP/IvEMy8dM8HcYbCcuGg8ecE2F2l1uRsNvy7KgU
97UFe83ybK0KM7klTd7FJXg7878OCdNA39qhTStI87flTpkr9607UR5VI3V1qRz7W7f4rFQhaa41
Bwtrhe2FmGojpsQyvnjwpHO0+BNolFbHXt9JbXguriyZix4WT9rmiH+6kLrC7o/WnXVPH2xPn9II
iWttOVfdq1/Ok+K95BymObGrmrGdf1FSV6Fdd/7F3ehtgOujHBJrElUuqFMDN3gtnM8JAiVk/7QJ
KR2yCwsXZf5UY5Ad/msZg97JK4gvXBNIuTgCtYYTc0A/duIVV0IdffKVn06xQiURZdDM+kuzxgX/
/G8Zgx/wcy7W2s5xPL4skWTn0uMeis7NzMj/r4FJ1JIeOpLhq85uoUnHmOn/A80GvTyFjSefkek6
sqEQ5xxN6I3bul836j+pueGGZWU8ukvZSbXN1SnmmKU8iebup8BEQ31s2Gz1vdE6LuEGyt0F5MmI
NyBJAS44iyHE3rYuCgFJPD6liTwCpbXUNf6ZbH/+f0drIROEb8xCSEgg1xjXgoZIdvdbWLDWf6Vj
AwyYQ0GyKq7aACMseG0luiyP5JzYGCgAEIPn7Xjv6mhwvfF2vX0VGt6HHS2ZJHvRFJw/UmFprxzq
esBKFRsSrDgKIQkzVqjRMOr2cRLK1vBqNOzdRnJaOqI8ORgdU2xsxeaG0c0BVQLc3+ttgRoQ0NEE
8iztcMBq0kQKptSByZretUBtFdeIXGAzDtb+aR/yhDEhCIEdQyS87GXyAvXciqfvV4QnmrLvpurF
rolEkb2FLZJxzNBUI5FKGdByi14YPeBowxU612Pm8Dyxf1/EcySkMg8cCvAmFws9tddU8WaNfgEj
NQKxWhdWHEzVRt9JJfhk0cfu5AJ5/q85kShlpULWjDxfMrkesu1kx5hQjZHFGCUpAujPUctMyKkh
BSmcQVGfUK/o+diRpfLSs3ky+3R7FWym/QQH5hPTP5FwxEDFW42+gP+VbR1+Cs4UrOYQZdzbtpq4
RVW62lQCukPrjZCzZ18W3p3mqMMi+gU6kdE2CGbbqPnUWuPBRsrWT8K8CPcFh8st28FW4e2WNYQR
UbUiJfLfQCc4jeZQ795L9UpgKNSxyiuU46d94pqHJPP0V1+xeYLd3PxTPfaKif2zDb3nphZnvv7B
PDU9FgYyBtTPNoENN6Jj1bHH3OxXI1Xss2iF3A1pg+CefqjxYxlFEtChuX0bKyzH6QHdz5F5YbtR
J/bprAPmtX7eo04ejd8cUKDL0NjWrtUcf8dVBJ8XXRWK/IMEsWzGXEPYXFCJZPlBP3v/9RWEHOle
+sVFtZI4pAFg3xuLbXpSPiNv//LBX2XpBuaeEY4/ZXKEcZ40J+EOs/Iu6MC1UukxabEbikQsCJBV
FoOtvLGSbIjOhHMZ36nE2pu3dOLAA1y07imkWUj+J0R/tNNSYsslk3Opdx/O6Wxfww6A3wJl3i79
8dnQHzv5LvmDfNc8Dcwt4YoHMRzRB13Ot+02zbxbEO7n8tQg2SfJZ+ljStMGFtWSd/QJyu3lHPnQ
MWb1WuWQv4cDsplDJb8QoXN6pLazzSoUD4kaYmDwcWg5YEW8bP0EwCZ/hB3XS7cPxG88y1q2R4cW
fv/Y0UmdywGrJzI2xV1puLvmzhr6Jzoz6Xel3LHQH/rEUdTXpIVy+LG0083SAohDjwWq02Wclo1W
uH/tEeu2kjPAyWZc2NiaTXEvU6e4OZ7z4FPvQdH3osQsr0ZXfoD9n5Tc28vstIq929gpBWFiQW4s
U7uJlDRW6er92ShCA6TtpsmvpVq9lj6Jjp8hbZuwayqTyt93sqDRem9hWPaXZkB7unt38xLyHqFj
w4FnKTJeuuMF3GhQz952KWbVKocYG7T92ej4F60CDkKT1OMQmJBqTvmcmgGjM+f6QXwMbhd1bLuX
e6swLNQnjcojDW7ifYIBElgYEKA8bA2VLP7PlEpLk5EV0kHm4mnaQi7GfAdL2idEqvSTM92Eiioa
C//9G0vderINK+JCnS5V0JrRRvOWzJBj7fM9mKxqdLPULRbtXST9swoeLutLyHfOQ7HeBpjJvCZF
yqy7kwX2cOu/ELES+LjeBAP2/oa/1XhspIgrNvZExkg+wbtMJ6l/vGaMsBT9YvJDFw5oG7ar+Uvb
NDmuqwdoytz1cXo0/FSQa4dAtfEfealWE1zkH5FnljUKfa+I0Z3Lt93hOj6z1vYBZuHH2kepDzSF
TVrGwtVpPhO+pWeIYiHAhXbfaw5I/Iu1WpFIp1UvxUin8YZgp945UEiR6+xFXi14e5bBLSkRhfKh
rbXYkP5s43tZRM+B1tTYZuD5+kAs8WiqRzvF3U5IFuZLg/Pk9n7SDL7AVQRrDtR0BOzGU47ZFDz+
+SDZQZT5UasLKniAzA0RcI8iOl8EMngABToP/AwK6nSpCRXi/o88UqTNqNFh+hNI1sKFDoIKOIWw
Ou4W8Tt5IOI+rWYly8pIGIkCy+B2b74/p9MReNyrpPBHWL6hrE+gsSRkwYBlUs7Mxo+wE6fs0Afi
jNsTQBkWd09xv/ud7Yd8kA97YJp/oRgRNKIe5LHpZd/yelKw9YDudStKpgkuA58KucUYbTW8+6yi
AKY85miUgTuIPWxF/gMD6rGOmoQEaCf2t5iK6r4hthEOQatMxsq8PFv4IYiV/MDCNxC4t84aJCO/
EqnrOTfgKLscS3/O9Zve8+gl3fBBbgad1yjFkks8gBFfg4v+LmSNA37EzDHW2fnsjPbINRvuTPcG
D3p90Nn0WM9J3FRumeLDv4Lyja7uyewsW4Wx0N9gupXP0sKMrZ+/v8UjyvJ86LP91zzw5pWSWYRh
xa+eJajSJHQUlBk5pLRHhf9VmLJlevLD7+8FVwFlNIv/vkVcO0Xxk/pqzsApc9zREAJr1H1MQ+iP
inEo9PKHj6HvZ0hzonN/Xxl3yMfhQQN7ak06xpS2LVuL2liLGA9NpiKH50/sDuxT3Se9Igcl8RnW
LmcYjIpl+D8TyMKbIKw3wyxWXk5sqw+vkvKkiyc6W6+8Xa0Ykdauvb2cb1DRzJ0UGSi+xzeg6Fn9
/lA1Q1prsxbJ6Sk+gRCHtWTt6MeAIMArbRjIspXlR1MhiSkSyhLp6bEvd8k7D1Zp2/fJBYiTuXgQ
jskYCdfJ+LlNo3dUsOTqfuf83YEGY+bdC/Wk/mEbRFcGERtZfJm90ZRo7/qcHZzrdDUZX5QOqLu6
F4LFNja72Q9Slda+LrfpBHbDoPli9XZ3EgGM4rD1n2DuZmVcK0VS0QeL84UgtLfAJhS4x9A6oOIb
6Pqe0rymXZmr92FxIWaonFN51afg05GTA0btoBburvxFGNDcOzBe5KnWyjaque/wA7BSUxOR/3De
vNx80BcKsHWzDYGz2Ao+hcSyD8By9FtPqFJjSjTUsVtQAHm8bui+ocQ+Up55BVXNwry3sDBd9qp+
l4piJ5gqoZyK3hxrhfn6fQrxWCLMPLj1wu1HPxEYMX9yDmTETpbmtksaK/HiKDF04P68LmvUnsvs
JCaI3iYVbfJUW4ZnVoCJWuGCwRtP/KZnEnTAplEtPy2ATqzaYa4SbOGBb+HM8x0Dpz0QQrlAXYay
EesDoDmbVNGKd6n7cOSPCM2W0+pFI6sY215ZWyTNaA6uK43tY9uwG5y1/Qw/hfrmdj5P8bVU1i6D
opJVgwS3J/YI9dEyOYuEl//CxN2yalA474575Vlyj5Ni6W3O5kPgfa7LN459bf7T4WLaX4VzdTeJ
NjTnBM9GdsNbfjsoWszHHftDSEJKxF7NfGGTuCKvsOyJZ/y8E7MZAo9jaOsN3EU6biOUKT61cU+m
lYDl2AVbccVQ69zUXpRum0+2mR1HVcmYwoWkWDU3ne52SKSblaUXG1wB7H3MktJnEwdEokR346fv
YELz6Y1g/tUPwtwpQk3pUrvW5Ym5vhvhjiasPoX6LwOwYFzioI1xnZteEpbwrMp4A85RJF9p+xtT
YGRwDXIoKecJatRpvHd0YDEtqb8db/JsPLKeEqSJgA2zwHOj+EMs/gZYWp+BSm+v9cKanN2w+nLn
ifkGMTe5aNRzp9vAI7xVMuHrhMBPr1THcsczoU1qoyU03oAG5ydgVkX5Drlvp198uTL2/njqfAWD
iGaapTSORblWj51toWksgT1vaXa8zaPT5tmrYztFwR0KFOfE5eiX84/wM6bk4AYgX5WlNVI1h7St
WJYo0/Xd5X0zAejSeYjUs8DuTHr52WPoXE5VaGpQ7TPWSguSxhamSzqAM+1Kdv1oBFKsMEBiC/c4
8s0mFvZz6ETFqx3yhTfljaNChXaMQTTwz20qe1BOTAz6RISBVIVWnWzFhmU8YgCACySnMazPEIuK
8HHhZv2ewsAAo6ErohVl3yDwLjVe71ZWxIcqlObd2vjXLrOYwBOIMw+Nn2qF218qQBd1Kz4+7LAR
imK20jW+RNPCANP2XUcVevBi7eRcZExEjRWzQqgREdrYZuS37p8jNbZVO3HW8yeR1fpM714vU1jo
Rdc8EBpkHg4quSpprVvedRpvfTiiWxNsPCAaELScRen69mbWiboNXAd6saZOD8T6Wp2T2vQdUXia
wKIVHdG6SYLrc2y1nGNOaSOC3AVmruplJ5k9K8LYfRaWlNoMYxGFjN/8Pwq+GbWBFjiKvsv8udAS
akW5X2YavMZTsH1vHuUMJkElhpVoKdS3hsWxLXQ6gqv7tD925sS4+c08hTrBe129PrVdPdOuYnc/
9wMGyc4lhz8LoqMCm99muMO7TJa3lO4GyuPcyDpTiXQZHRJu30N4YpYXqk7ren7BYUhAhjfelZ7z
g7TJyLT/UnB+ryZ5aUvUas8TtbXOpfJ4vSZYZ1U2YFE9JouRcCE8nRl94Ke8sUTIXoQuGGzuleQB
rr9OPltfZ5g3fxXRefak6j3YkvJ+SQW5J51qE98+MCuUGM2q7PhdXBqik5AHnTVGz/yoS7mKxjLV
gzgRxmmYUpEziyKrvDgURajgdVNBhq8PuooTDh7zzmPlyDy5miNczgcHY+wzUr53LDmFJLSemdGi
FDNNa58Xy2CWmQm0x0gmeiMm4bPJ9sGDYvRndhapyKiIsO0F161B4lZwm2S1Jh232BpGTy3eYKfV
wNgOKmso/x52m5PALie+vByQ9+L739Q4RRs4fDDfPy/Fv/uJevSmiGryLkMasI49+5iBbZ6HvzpK
xkoDf6XE0evFnGO+ylU5WbrAy5qwaO0X62LyhXfc+ti7d0pp1LvsrYm4b6naIXwSGqSeCGuv/1Zt
F8PKX1GBhHQO1XrN0zvlWsmXY5iunJ54b0tw7oP1UB+jszizuFK+HAwg68ia0BgmpgPQOFeiEPlr
inI4YPeccxYPxe6XTyxmeUjLUtoivvq0dnjmLx5iMhfbslf11mB3hlaRv9dS39DDVpb2wC0TxS90
UhBGHtN3MRQAhY7nXAqIDZuK8414t0cfz9OZNxNxJcb/xqs/933VkhwqprWkcl7XdWbKmPU6sBkl
9xZVmU1WSVdFgaI6BcunvZfDGBxzfw2XMDxTUOKKf4qfYfFe2hzdnCeQeZbY5AEUE50Y+Q62GDV5
r6XRN/OE5htHGhUFCw5JY+HgZ+0HCi8ltbFEMgSRQ6HELqGFsJ1KBp3cRg8ZUTYP90RNhJf0Aydq
wdBVT77HQfe8NZfgAiZ28qe8TVG74DsGT0gp8QH4+qCWNb6ehwPscEkK95RpV+n8bf5XRlGg05G7
qjOxr7jbHavmoeum3xBJ/BpgVrk6CzBvMUN2E4mqpcCjmC7DTynKvd66qYEom1NjrDcebvcMfTyo
fsKSTljAZIwfWiS5RiB70GxhTXkjD13p/OrAXznhdeBffNoGOfWOCCSqGbITLPykEYNEZks/xKrH
SJ6ers4ZoNG9yTNnn1pPWQjCZlQLfUcxS+fGt7vkW+L5oBhvoqhJMf6dRohWJ28ua0CFFkU1psLQ
KOrN799gSY0deCw3Fb9wEf3gF8991uul2jKmcImwNwzPszb0CzFN3am3CnO/MJZSmrbTt4D8XIXr
BmXFwjF+Z3IQY3vodnMXh+v60HusOKfdqOpsOSSYQtyUNHlFbejlYTbAFa9rrtqDCwjeV4e8A+nx
qyg29crCFl9CtVUx06bIY6DCG6JY06wa+btpuXc5aclzFqyi/QSURsG1RyOhMw9P6b+Su0Y0SmZ9
sYZWeBU1bHtiYweMHDWE6di3iB7NfJCubqtBhoPK3GkJuD+7F7spb8JFEJlTabAEQCSc+fW5ZfyH
MG0nzuDzcWiO+5Mtv3r7WnpboC8xEveOUSJ4MLbrec0JBCVT+ayUTNEB1Zy2MTayur+HRb52AQIP
q6HXMCeQCxxlveO4QvYJG5mO1651qFsCfAcjTDT4BebeCchzHiJLapdkuC2q0MCqLSbNHpBH09SI
kN7rFDmBPc1fU8idbD8ePgMw/ajtLr9CGGzwpJ0fkJci8MMfeDo/CF9mCHTZJhsVERmsDvhFxztJ
0ot7lWwxn+fHtWOfqk/Ax8eLGLtZ+sQQMDq6i7HgTvUfcrNCB+RQhFXfJ7RSt2CP727A5RKTRbjL
sLliTcsDWOGVYkyo7DQnnV34fl+RSPIeYCco22Bhr8wUK9tZ1RA4pGP5NOxuWAdXvEW+vFBDvgrA
CLnL/sCr/Rc4FcdcOJNlFNwc0mZIyF4aHN09YMlN0lU9zNEAzWmgE3BA5oIA1Fd80Z4efdpNIAEq
yoY8OJRhgT9G8sNva9wNBbm/5MiHUUO6G3KfjgaDGLzN/H5TzgnXcNhHjK8nyzfJ8lAzLaOx16wj
gS7G0W1XYnGgFFkkhpqgZ3GAxe3ye8/CKUQMAaXw+PsDsGsryzUJHnTJCe1udhqTEFRi5tQskkDO
gwEY8/5cftncWUQdaGeNTDvxO5sAxp7vRoesIpnl5D8FPBLyEa0Yv2UaJ9/Aw/Zp9SAUAY2D87hQ
f78RZEdU8E3BMKq0LwezlnqekodhhDAGUt9ymvrAksCfiYBIXMTSdVQSKQ1UE6vsRA7uT9NZLTKi
6j/hjGtGX5TFkA4xKrdqOfYiH7EkjMi0Tr8kGdHuCq/NW7O7rWcU2VDWsQxvpBxMBMu5myssLCeN
fj0Jft/AztDTob7H+8Qrf0N/Z+sx73TkKtFL35vKh96OACG12bTZ30RPAwjUmIQi/pEoudnakL3y
6miOlsfSQKg5mYH3K/2VorWokwpgcwgMq6G+OvbF1Csq2Fbj+S8sWEOJ20vclTILTr7pLNd+YZJ+
7oL+dlR9QiHg2pXHz72NI18jc7VofM4DWDS418OLisLSNkJLBUM/lYt/yy4YyKCtXKBpNcdyNh6p
B9rrMQ1l51RPx3FcdjHKhOuI2pwAiS++iSvJrtDO8RBEQpyfzqLEgoE+ASVr3thMJKEmeUtFEDA0
Qhchn9gg0MKJ9526yrhAsDrA88HHLIB65ejqyxmgo9WMl6ymi8FFdFoLvW3W6h5qx/sp08Ud4TQP
Wfl9cBh/Vqh85fEqRMBnHPb82Io08MB4UHzSXeBkbZXBNe3uKLWYQGKDZBtlrnLW7M1hcyf4CaEf
sYIYx1VIL4iHZ2rnp/DWNzJxMB30A6UDn/rp5oFyugFspxdFCi+ozChTaROmXv5lUWsRUQu3WHmF
bHmy1xW/ovpa4u9T9cgfbhBm8Nus+RdfglztOPC0J8hrZ+j3lwygHecqolan6V7oqt+msI2M0MCD
PRVxFZsSuQ7UrVgo0uzLrMf2+DgYO6j9txCAzfmJT2qW0YCHCtEEPY8RNe+W+rQtvETwopo1PHth
/UTmi+pYNlhbABbRqJSGjZsI41D9Toklm7YT37BieOxIKpsuDzD5h+oEw9V0h/aOLr5UaB6S3Z3w
I2r+mwwU1IG2uwvEXmPDW6IkqUteMgsINyswKp68nw0qa+fEPOpDgivoPeS9CV16vKDYMKKHSySC
Enge58x9jDT0FHk+EwZSBKv+VbK7jgEWgWGPXCSkzEN7LNUX+piJyGOQjd41g9YC4xTBI5YIGp7i
6clUoat9nn6P5SKIyKa+mCWfH9lBZ6iFdg9a16DKAiRMBNKatnPdVf88CT5zOFHdbvUew37BiWBS
rTtSH8MtQDbRTEg37rrZpZu8/omhNDgiFAYhsN0YNGmCoAfAYoZoHj5loOUpnG1WSBhCQapG3c9f
Dy/VMlbzDZLEfPEzz20ETxNO2WUtAAjuRaAeuMY9f8SxirKwDLwmHOtMEGPCBi/V9HvQrpf5dUnl
Nyv+2BKMbQTXlnSJQquXE6h4UnKnbD8SfKzi8Rv9jywq4ltchSDmLd8O1B5Lguyv6XfQ1QiOWzSp
0dRHrldDnTYUxAgX6NaEMs6d05DLI//1bksp8p2NBPTejnThCGL96lbfaX9OyHb3YcypGA4y7Ob5
Z88RdHIKe/L9p43TCdretFaYwqw3uirlBSLBo29gltw3dx3V0uIjPv+6zjpHxnLw+0EorhQ3jxLT
s1RZu85mSLoMJ9fosKs0BshdUNxv7nCigOXZkXqdKEyvwuS8XO/NjYJL/frm6YwQwe41BjlhnFVJ
WSmVtxpufpb7t/DaVfTZZ0TP7wDnYEahOeaEGUiFY9383OBh9akA/0OV7daNAeCJfkVkbI2cOH0G
owvb4NrBWsHqiWB4inKMxwGmU/a7w4blAdbPHtpsjcbFNmfKZkt0ry8iA5IPlFeITL6OyQMQwbsC
jCwkaKqUS8tH7QYtdpDgP5HBLepHeyg5ekigaE6Vlap/ZerUf3kjIJU9UA0ukQH4oBmDkR6oAkyb
4Jfcnh4COJ8xm0q2YFmYUWeUM4oas/NPxWLIOvLiPthG3ZmZgOaMhN+2QZcoYrIOtZvX7fnpysTT
uAdws2IvSrOgIhD0G+XsnwL07k7oOGLnZ+Fc5NUfmXURHe4tz/IT2jAg3uaqpW+V8k+XnTrcsFrg
7JJU1naIa6Hl2jFXvjZYCSEsVu3bGqG3n9jY2D3G9Z7v6kGUoetRKjqYgNLJqli6Y7DOrhrBb4dT
DKaffS31BbXRS4h26jKnzj0E6EXjDA3miDHLDtgOz3ZWRgulya4phq8vzaLU0jom8PD9+PeTI0vD
l5cXdx0/cmaJHWkF5mFbPkFQd121VxA8My2XO570eM+ezE9cT2B1BSSbm7YBXAbk4DGy0yD3C4m1
pnXuk23ToSBnwh+z6q8j8XxPyC+Qt16cHPu28CIsbnYM6yE6543wxGlTBjLmniYmCh4ZSzHHhgs6
FlrHX95Lmr7sxVNwbUAP6+8yqKxN2O6EocFRoJcGcy6r684eukjBODW2hHroyy0MtqWvOuaWJZOs
gRXsXkwMzW18tO+13CRTuEp+M4oXuHN/4B7PEjV8DuGn1X6cjchvr1tl2+iePBPQ85mwYCq0sYrY
guIMREOe7/zXhStQrDlSad4/3cuFCWt/Ix/2F12748GDdYSon+IAZ6UOYdYtPEneV//0ywXoMQFA
E++7+wS1F+3OM12T5TgLjfDtQYMaJ7iwJkK4NBMffhtfuxRmIjHaBiGTTWEAbiBFE7YQd8Zkh/i+
nRsUHHdejotBh7L9HJF1I9Ddx4uip88FpQ4P3A+C+z2b4/DhQBGNpYkkHdUDwhdI3Aq0zim8Pfgs
a6wZsqCR6WU6UB+6tS46g3tyLG1fncKN10wy3+ajFoZrrK2yMCDbnU2bpwrFgmE90IfE0dRGeK5A
Thcr5M+1mFwDfFKY9Du4HiDPtt/jn6FDSDYOnB1aEwNlaa6fDJIENfI1x2VsncHja8pWSYpMrzvJ
Z30kqf1p9AqAeKCFw4sV7lLWinkk0rkAtgdOKpRg7gcXGN2RNYnbZqYZFs9AGCgYVRsfTL7FX97I
StsLJAMotFCneE9Y5WwW2ZN8obMHXkyZgrNHaJidHMBEObqq3OtSOC0I3fX0k3ClzpFeETppJcrP
WsiZXWzh7t5G9iI03WIU9xUirOlS4ko8seCp3IBqXrB/wwxff1AoSUeSVohaYO0gU1UUoCuAv5Hm
jOQv4lJpwgsEUBAC01OISmQJAnNkJGBAkCY2jOWRB0UA9C05puDUbj+xl93khnot6xNGcuqmAPDB
7iKafma30yXmnw+FQrMGxI9I6TWiNfx36VbxebiGvlMC2mHs3hMS1f+3N7MJfRBzFsmqWxeu8Sk9
EpW88Okjck6HShrDueqDAwVp4DPQgZu8R9EELw57nXRN4dBVNmYfZSyFhgzCGSCuankqo38Il7LX
1xwbFLdRxErcaLK71CBXGCbQ7eEyXixp/2miIAKEw/wQMEahdk1MwFwANCBNQIskKGmxA+CSSzI1
NBq4A9yBF4VkkcK2jwtO16IyAiFR8nKHOKeU34+dsgYKSc/SJAK1aTpWe6e9PubIWAkWPTwpBW65
RRmBY8KGggR2vUi2CBNdZy5XsCeRv5W1bpSzCIGI0PALN0Q50nuoRaXq1eKiVAUBvXKnXF9pX9AZ
A/zLT1i4r/KxFXCaB5BcFDY8VWCqGNogt+lzicVnRwryt5NwcjSMTd48qrwOjKe74itxxt0ZxixD
5dKQDKnRTfGZ5FyF4sYy6aXLJSpzm2BZw2zFYQERhYZNenlPQtdWZIKhbQhBnPrxUAPXOEm9+VSE
lwdZ3IfeEL9jJFzGOdbcSHOQAhPLOuzl8ERrbu3OjbEaqajUBSRARF/DpGE8B5d3iDBHD1KQtbvF
tdfGYoSLHdmEMIX6aIN3Syiv5TDo43Knn6ma/jCXiDmiNz+Q6Moawnhev621Iw5D/4wiHyBm/7ih
kWs6l5jE1DjO03EJBT18/t4VCbCr4ySzznXjHqPkjtklGEnWvZd6iK/9MI9ex4y0O0rj2QpCG9wy
WTOoP/GOumONsfZtCn5Fqhp0yNQ8Q5rIuxA9sTmShRj/t1ikBfN8fcNU1g5zLDBzG1LWlXiOeiZw
HnzqRcB12osWn3GwNvv3aff5+Xi66pB+ComMgCbAsdKfJ20afEe2qzo0fS6QPDzCZSVoKQC4hqdY
JRCTBsUoMRcaBuC102VClBezOrvfuNLTFhStJyMFsVk0odzeeVsCMt/Nsp9sjIfYsoisTIF18Ouh
G51bmKF5d0CK1s0yjwQiexaFAn3huXRXW+mhf232/NRkhrooxXaHTbRqo5Y2vsW7/7UuZQDAOB2F
F1mb9hOhdX6SAyCdaMvIAnHW5RiuRMYaK3vkyjBT4Ea1Bb8tQu0IYew6v/gYFSPkuHzfItHxoAti
3zLTlOmN0QkpOaYmcj1641P4abseZmJplAWdqx9Y1D19mxb4Wx+ZZYZrpSvCQHpqwihFrdd0p6r0
mc/Va0FidkGTFxBn5DuOLU/AGXPx9psvTmNpOpH13UM6QINZBdE8UPSpMoiRt++P0bvd+ko9MF4m
XueA5yuKbrduLQYa78kVFIT9g7NK925eWhywJToYA+kwyarWZtMXTnKZjScvTGDtyf4Fjtr3CZ0w
5AV0FzZFH2Uty5AJ+pH92ZV7zlyrWTvW41TpBfh8waQzGjKBVgO1lsZmzw3up02QMYENL5MYkk+V
Yj0qePWHyL8vqkEai6lLukhL8RzdDiRQjGwdCSKPZ5ZXuonNynVwLSOdF7gT6CPvZQr8tzSPdZye
2SddhBe329ivHNBF/26QkxKLaSfZdhRNLq3UDo4emv1scRZQU82T7vE9rUskd3EtVArSDag5Jjud
QOpuMiMu310JzNuDiZom61BmIwEKx1JOI8+y49yuyAnX3NKRS7pYHkkasDN9x/3uCABLXcYMWSt2
XvqkJ+zkCDFnCzoE8IsoklYwHRhAZ7RrKNHQZlx2oIbd66UZtUWZwIRFjubkJ5ZmhgBypTAAS0b0
LQuEDa0wTjFmcxST3iSq7j1pRmBlf2RZWbUGMiBrIAXZM36RZfFMocTdsavde91NlYjEeZ8y+eid
kpe6swE6+Mlryhlh4ivgQxRm/BUMqvYd0K9kB/6zY0vMY4nSzUZnkNCqdZOm+d513pudAsHBP9Dk
VfjMv9Do6oU4ksmtK8IaoKdgPotAjAaRtvEx7c5zgSLERnNLyhcOT5eVc4vfxLGGwQb2H6yOYIQO
zB5m5tBJYqkqBsrmfpTvE6TnnoN49vMX6DfixeudXtc9vDFTJwSDdP4AGDFkebLWpHm7ncb4xN6S
QUD8KdIkuV9fgQlybK3tkU809CoZXtMqBxmYE2MnOgbkSKBnbDBSdfW9OnZIcKDj97yLMCKzwkZA
iGgp4SaqUbqKVE8/yeDb54UY7UOFCzSPzBhQcXp36iZUg24G1w/dm0WIB04XIQq4gnQF71rBbvVf
lhs/LkvGUv6lvYJLXbwLXN7n9gV+DTCuOaypzByymf/ume7ULG8Utjs8kaAEHnNAOP5L/tHjar8T
i3MyJm8EwQ7tduLo5T/i3qlgP7QA29nQ3J1/tCHddQQ7WuayvZ23ueQ+oFf8Bk95DZubdH4OHzSG
5i/X+tzioStAiBuua4qjxZOcOwPtLxj+6zPlFYJ0ReSEcl+iqKYRrVeXul4qa0RH2NGDsBXkWU2f
AWfXWn2aDNK1jg6Isuz+mEfYqUIQZD770GJVCkWSaBp0XGlL3pYyu86DMkyDM1B0tNX4BuuR6MJi
PCkL6Jjm0o9K0xTBId1MO2QjomIyLmAlWdp8s9n5bu+RLFGnH9QwFX7WsWbcPWO+yI14/AoOyjK0
PyTazwTte9o0EOgWjydKdHx/218HgIqiXCF0Ofm6U4D0t0Hnl4xyjZwOgKP7b0mAnKqAgQxXR+X4
+UE+SE+yMVpU4YhLzcXH5+ONcgYcjGWPoqNpbanFwijfi4X+USJLGjn/+px3/4+OKoretsDWIJqp
DG/HfS3PCtLH7QLlOpRjnPGN+M/NoQ65dYZeq8Gwd37BD+7JWFbltu1CVhhE94QpjjVMY/FwUc/y
p1u+kgMegkH4LqQ+ydQ4+7VVsji/BzHmsmdTFbBsOD6s5JqjWcN5OYx6MtFwdRMiEVfMgfFhN4J2
HlgbdBwNVzNn5sEve/WHIeITx09d/tlrKfozYevi9EfL2cJSZQcGa6jcmXnZ9Gs5IPLfM5N0akvN
olIlIEty218UccpbKPephmZU9U6mn+eZwcXWludLdn1qUS4fh1l9TuaYzj8XIGy1HMvuqR80oF6X
V7PBobSyVDjXaxPGRObL/6oadcuqHn40CbgIS84OR/paooIMqSroWwBwIH2KMsFkW45o8K8MVrUo
yzscjnhw++zRVfqE/yJxlFentWz9sZKQ110Z1lt+ueGmVpe/LBPfho/i9b6r2fwymOVTIipBpcvl
SoWagI/seP8f18Y5UMamY3AHSW7S6TQ2dlLBf2LmBGFwVCwbbFuU9dPb/n6CTvXPDCmvGW8is1D9
D3jSjK4bOVsKh7XR/AuS1bTziZMXO4bjPl2JChUxDtA3d+3c4mcBYDy2u7DzWXoC7HJ9sin+43ep
XUsvDzUQc5nPynq4fOB5f6W3ajBDLNYGzcfd7XdLA+U/sODazBddFtCQaSWB3nWovbF4uGVGX1HZ
+GgfUXVIbLtQte2ms+FfEN+mKGhj6MOczYIO626zs4cflaK1rMRoaE7DLYxLpctYYSr6R2roBOTE
GbgiP/l1Iag3WvdA87ozrYeW5v43xQQAxWjzXfFF40loREKepCc7waY1v7nDNJCcJxpMulKXkN1A
74/Nc+D6SoTZJoXD3L0LwEqobUes+/XjAjV4EdzusLK/e9fZhI+NZs94GDVr/pWSi/Ibo336CtS9
V2v96l1Mosjgo3+9H9C0qQTxmYMRPC06WLlAvoe+6b+XA0L7m8tUfRvpGBkZ11IwzoUxOLget1ed
37Fy8NXZtH8c5P1onGt7JpMXS+VJl/TAlM709JUs2FfI+Yymh6Ohc2bcaWXHp9Ywh/wh5oMkRzzO
Mp99lR5LZSpwQsjyzntR1whEqIR22bN6giNhKYanbxxTs/SjX2pO3CvebaNu3nlBohg3GfBuv/rm
vxt+br+22ErakKVTPdbYwT7ds36B0D7eMM9c65WchTIcUKqXOG0bhFoyD4WFtsxFsecRC8iIhNbN
NdXK6PHRWmQoxafojT+pWcnM51AjjMHXJan5iqhUVHACPQN1I5lQveLt8yDZDHty9Ogs75u7AX8x
au8Ni2WdJMVjhCC+qxHId7OO74wld7nDEu7n7IsPgrsbkX1mdel3qQXc8Wj849qG/GrRolDFV+db
expRUuqUXBf/l9nqLl8JEoPvaUUPTUYn14OwT9GMgY9icA2hGolN0YpWwddUzmgUdB86cv1ofnuf
tv87yxqn3TeSRtQynDONs589G2z0zHOScmVe6mbXbxDqjlgcmZ0rZst5Mkr7oyaHJMCoYywvxpvk
MYlLJ3GHFcoy31LDn1pSnYYnn1bAhqVtuvk3qmX3D5XmzpUQ21GjD1Xsf+fnROMRZiGF6x5Ropoh
aQXFRj/YG85bH89yM8gXs9+L+W58eu5Aj2iQM7Y8YXaLvRYJ08XZsP5H6MhKG/j1R13rmKTi2zyl
tmvL519OYb2UBVapD/9BqxxjV1w0JgOQShMmSL45PCHiqVEFJpt3HXrp9338HRuFHCcbdqVOxrGD
7px2uueF4N0DDol9MNGXa4kiZjOcxsG1xks1YM+py6jy2GUfUAQSQpUom0H/cfPjnkr1b47ThI2U
y6nxNShEeB9laMA4tx3JtiDzDt6pUMIt5WwjqbZnCAANh6weODS0fZHwFCmptiyWa5wfBJsG3kri
pkzrwUs9zIPiNH8LX2ZOlc07Qknp7ZitxpWO1EOkjMqZwPDhgHSGOPpznTC8tOxnjjCPQdiFTDkS
BfPQkcMxgulZJMPxVKNvqyFwX5Kwr18ilQsVhlQAa+rgPDmPpEDP0POJxLh1mtw/FHXheiQHcy0+
GPBvNhWiXZXx27PbOXxuz1uKb8oosotuu1FSBjXp8KW6NHO9q8rGO1CGzvhWZ9ZomAx1hU9wVSWU
IJ+S+qs8iHGMfGhlWn5cbgpD0RoqZm2Zscxi/4EddegwRY2xd8R7MveNnd+sAK/dlX/p/ZmLiPJ+
0N0Epd96m9Sx5In6lkJ+5VY+d5rsLMkcJMZUchGRinNppCWZWre6Sfz4s/vRalUKqd0cJCKamm4n
vmfSgceVEcLcAXzWk4uJZ+P7oSnwq/tLNcHW7CKtwc1zm+PJyTYOHzcryOHIYbgKNXmwTidXBjOr
coBzX9eo/0KAKzbmKaQdlaRwyq6PQdLwVZgBUV6ObPGlQ0Xrz8mCPNQYXpBs85xWV3ojQpwc4gqs
zuY2C98XH27N8oWCwkn1JX8UcyK5IaByI6KCT1QtAqkxAjiToPSi5jUrP2R86EfBgqsijQtMJyjP
lQCXSsxurO0XLPyHVsPcYShJujNArNsdEDw88SL6ze3EKY23i+qgSO9fdHZ2WgxILCur2UB5fiu0
9thZW1VVXv/7TDHlp7jCQhzz/QHZhFZEyVkaNoo7paHtgEQgW2HWv9Cw66G7Rw64D26sCDRoTGuY
aHOygE7pWJO92arXfJZ5hvdt3pqod/qbyH1QwfEWcpGVuNKP9NxGhABXtYx3PUPo53hDNfy+kUMO
3zMO/G0cyYw9LJCHo8sSKBV6rsNbqDeJu6kGLrXGYROGd7CmdDXaS2NOt47Sse1716WqZKVyIISh
KnKQ9vr3Wuk/JD64cSIOItkUEgt8+wH+7qORkCeeC3eotSjERNzae8XTNZ7fRcjid3d5UaoS2gW8
BXziKY6WiWSNbDGF79FyJOuKCMdvak9hgZ/sCTPRGUYmzqoWvKQxx88cKM8KBoBTihjfn71U3Vj1
0p1zzbuBp3qId6OoKtZgRgELNHNH2qMAjJ/vwgUjYhyqaVWi/1sCjlLoo48j0AuMaqguXs3rKppE
GpBHFAmNtjAm596bxroffDRK+2hIhgNeY/X1X45fjy7rCC17SYpcWTeoEbqw3dEI7wpDfA4JiQ3n
wNzAHXf+LWepXCVjha6QPcoqGqoDV2C1P4WRap1A2+y19SBwbZwZdGRY6tqQVtCNt7iYXdMHDUf0
TTXrSSYNndtSPrkjvz68APe/9FMFGLb5VokAWyUsxr/pDXBHQL+zAfdPWJ4BuQswfk006KBE48gJ
MxKOx4NbegtjLSBJpLJo7Pk3uBN3y4Un9O2fCfm0ritIgpuCq5XVuWXPD+551WyNilRUV95I9TuA
R673muq8vIVPjed68qPi2p0FjO+OyojiCNrw1Di1WYXdmgxIFn1L/znQUDV7XHeoR92VKHhoMxMO
iWRe7Lh1elzkcIcLGCHVB17f5PWcB3vhZYcoY6GBAqns3AKk5T0BdNOQ4KzZ3rQoHUGs5P9XvAYX
i3u8VU++v3k15JYQlau8+FviSVaQl7aVo8rXpKhS2hMdL0rRVCYW4psJWWuJj/sfXyp66k5JBtkC
X1W+GWQICRcBQavHIlzP/oL8R+FZoqoSACH1ZaUw/DE+OcIFexnUCl7j2d9cu7x0v45to0PPZiLy
dns1Pl94k8+lEnrQlmgy5UCazPpReUqpj4Sn5S/I6oqAGrT6rrCODpb4kvGsft3hL8kmJrfXWd2C
8Kuru+jTXRCMA6Gt4vIwQ8G0mzbjxW8TPo+S319rBVpk33Ys8IlB6T7fkSG4bTz2us//nlXbllwv
cNSyN29N4oTqPOhZ6YcEk3QnnX++l/cdcxZGewH0JAqojGSaJxYo8bumoKW/VQi1qy2aVRdB40BC
3qB7plb9tNYFZKZPNia9i5aSRO73+j9ChPSSMSufz/kkID0Is9U3ptxeCYUBG4xB8iwTvM7vZWs7
UamAjskSaKsUX1doCoatRsV9pkcuGPCEdT+PLFWUt1LSzcvjf9SWKoSX/ulcXNb9ZRMFDzbQWGJN
DaOuRMIjqFlIrRLpeEnj3lP90M+bxsV3KKOHfVPuwT8NCNv9+VB9/zmGSUIu+SA+MMyuNrm8s/Zx
c/iHvF7IM4GlU/Ao6UvVHPxqkNSRMqyPz89sUjF2CLJ8jsbdhccCq27IupDvNvKyqq8c2OitV3RV
QlFmcGoEHJnk4iZgyGobPBHlZ4UWoJ3+NBe3CldeigpoZmUpxQIYsNh1TkYNrMn+g/6jVxXnGUSs
slP0niMmHYq4yxlK6fNkFsLT7I8QKcjBZEEimlqjsq0DAhVjAZ3Z9AA0JCimCQhqjHnsEDurharY
YsePLDIen5ThtKrEi/fjGBnS7SPGIE6ILKAvu/9fMs5x+YQaFAaLWSIKJa8j5CQsq16+EKBIs1OK
q07Am83uapKGvP8YSimKXN+kKV8EQ3ILhHZtU3A8rDbjT2sZSEoWgAp9RQ0nRixAsjTj2XYlbGDF
woBqLqMfRVTpFNmPMffZHQ//H60zT2iIXJeDFQjjvswh80atFL7GNF9TzbGUwOenFLSKzI85vRHN
yZTwdrsfgmsX3snWfc81OJulc0PXia1cQxcmyuf1WJUjUVYYVuA1H6Mtv2VIktqFTcVAW4VNGki2
Qu4PMt1u7pPEpCTOAoNvLGJxL26ipRooKfI4DOSFjnu9iH6ydmY+s0UAWli5VJsXTPHWiH8iNCwT
e2Zau09E27ZHCUIvGg0LRLVVOHHl9tiGGBW0ILpXQNp50chng3bFlPeklE0Jp0/Pw5b8wIcWJOBO
SLtEsM9RfhgrvMuRX1Ivgqo/Q+DnnYrK/f4CY/Gfjj5ysX5K2Vrva70v0qtQbhUTbuXWVRpmoFyc
P2zNV5Aa+1HQQmtkeMAGSdrE9jOPXH173+g0CIqf+UPyHpWA494Q4cJWxPFs3UiOed3ejQWr55IN
jhRAmEjWrCpROfEIPP5EmyXdkNCsDIOnaNYDL/xE1nmCGVTf/M09jFr8q3FsQkz25N0gzlEkJ1CA
eHSRJgCAVEBCcwFkPVDjwcZncJeVXMuUOtOGpmIiGoD8fR7CGkG59R/FoxxteyBfR9cvwRdpLHU6
yEfclx/fDrTkq0xHwY3UOEhTB+xSHTbi3KDj79emIQ9i9X0Rj8jek+Y/H0SYuxffMy5aaq4ZpqZd
/KvZhBCu1TgJXyzZV/G6kwtEaNeCXyvJ4X254j7dLZgh5YNtl+9dW303Py46FM7rs5k71/aBvHhY
0BkM0KIO6+aeJecWdf9lXZMNT+tg87LA7g1boxydNLccxsGFFiStToiVT2Q9hh4GHgF1XWh8fg09
fgi0y4ZsxeOKFUZTMgDNwkcXicFS4gh3FVe+xZKnduzbONcIogLDb4Ra1z3BAA5PcAPJo6fWAEq5
uIEi7dtG+yDr5Gd5jXRsOud83bL2B8eSfeXeLDrD2QbcCCqI//ad0eJrOWZsliGLSNT9yKjNN+qJ
iMjqKNUaoDvSDP9LRqEQZBX2AiPl6Xo8hgFRTSEozf6meyaoxzmWPlv5Q36SwJI8zRy8GjVvmOQo
boOgAJtb5ck8ln25AeeBt5D3ApVXMx2HhJwTVgRG5DE6C7VtmNxWnGs19NX4Snp/s6T4huooG+qx
Nmm7JeEaWH+uqBruTDUisTIInIDlbkXuAmcHmnBeFwweqGZ0VKAn5TT+0NutLu+o3dsHNVLsvAJ+
7/4LRWFNO1DupfD4XHyCAth6ZNlDdvlQBFlzOIhNtU9m2+cOQyGNRox223pUy65dg7mRk/QbgvoU
RJkwCsTf4yUKgvE0yxCH5WPHuUjpQcq2alDJ87RTsiLMrUop31SeQTWX4+H6lMxhb7NMWJZQaoeC
YlM8leoAjiwsH7uzvwltEin8tmQIcwnRuewCzdLZVUcpr3nWNQ//gNRJVY8iWftgk+Dy1t4J6hRs
6P/X6D6x/m8P6PCg4Jyli3dXWlgK9+I9GIP1VJvkuvbMoT1Da1a1b8e8iiE37+AusFh704dxLnAZ
CKpNzA8zbTdkr+A32hgDZYtjHZOk6/qq36bT7ad6PYFQ4EcWmOaVjQD3EBJI9fwjPjaMHaRLrNXL
dcjqnygaYNxVC038da6iBR9HOo5lKFzmuR/vfBajQqWkVawX9UPf4bxc/AaX3KN0on2coP/2qF9c
N4LtNXEy5612xNBiehqX0cNgKZctM+269X0CifRwYRstogpZBxw19h+rhKhYNtN3O4iSS1QNSDrw
JODEhiNpIdds364WRWM3sZs97FCRGgksXsObKhsNZ7wLguPly+6BivNzEclYKF3qFUWWOfsTjf7G
JJbirSmkF1kbaHCuLc3tqCakoHX576zx29lS/10YBQk5dobOfAOqao9Ka6BLuNpp9aAOj2i99U3r
uDMocnyah+nZJ+ohAFD/WHRq2xSd/Jy3/HBJK0EcK5sQTbw4O8Bp8mhPTOltJAEE3aU7IKHvEiiO
oEoYJbhQBP0QSdg4gxtcxaB3hF09N5zcrIP2A8RpseEBzeshiBAswBmXb866zJysh87QvKgb/9VG
M6hCaQzXQQ6eACtIsGJcpK+CkYJFq9vCg+9RG+CWfDC2enK7mBZ+gBbv3TdlLWkP9Wq1REqoMnMV
5xi9ABApGui2oV1O5cJ2JMlm7fPd9et3x/nkkAkk5dsK/6rG5+gIalJX/9dkZ3fO8/5en+C9Hs8v
nVlKcByz4RmPjU9zSOpt/SrpwBatIdml7fXQChCO6jz1Lw7uBRX7c3fQ2xp4YZHTmzNw2uIz78WG
rmXnRyx+x0LWc03SsoaObN/02DMoaMgf2tDHbZWi6cnwRPguKgUu/KErDzCx/tbnjx7pW4JdGd5/
RBoswFK4U7OsX1btO1cY+RanaPAoMNFfUxO6Iig9lE58x0DX1hP0T8qRRtuxqWrxf+5+167LNaRG
MQviCzUMHQChW6IELN6KlZ3JbEAX3d6ACX5mWyyz4WI3tz6SqVMCx9qyF87xBSBT97dF2quY7lNu
YyosXDuEFOmhArXxEPGkh8awJOsbjIY7T+x8NETs5H5TEcPUaK8eLkP+O21QXIrYk3zQsRkF2f8e
vIV95hKN38Mh9uY+M2qMo41luGf0cboe9ylP0WJqVvBDYcp5Y0pKLGGs0yMsye8e7CJGyBwCMtLs
St6mOtSQZjxpiiGFM84CNaa7CQyT6uVewxw7HsHhzlJRgopuTiHRru3eW/vBn/ysOQi8EpK0+WrO
EFnQeKGr1elvxsQoypaXic6VQUGT79Xp3YKhwmisUhZ5+0RDVgn1wP7HjsWSxXmiHkb+k7DJxMhR
0/h5nSP+pxOQMofI5DNJiZZ/AAjy2di/lYbNPcqvLKyQyT0gKq2toI32kWDJwJZmMK7mOfuO2byK
kLYUb7vwJJg4xjiLXkbKCrKgVGbIc81yHsiu78dMZRALFRWFl1HrigF5Tu9UwXzXXShokwengsjU
mYhEnkvjTkGMC8ZnZ3evetwcq4eGEFfGWXVRbQ0N1zYEentSV8jvFlX0H9pZbtibfQYmchkO629E
jch8dNTwOn58XV3kJMxfkM5oY4gffGPTZj4ZTFikrbIaR94evLqU9XkHuHDDo9ZjIfic7OnFUf7t
AGjTfghUunQPRCdvMg7I0KX8UKIsLdyOvyFF31EWhLt+JBR64gQj5xgXdlqkvwadespWra3d6BYq
LQRcbv8p94/U/Nncg4F/g2ryMc7gYY38onaCCfyjiPqncX0auqW7WUfp6qvMCT54j6yzzScDWxAI
2uxHKFWSYKdNa23bayOK/1vhRiSBr/jD1aZDNT+ekFhAHjJ/pd1CygHUKh/NNsbZi0XqEYSdw+vb
Cd56lomW/Ki0t09i4tLFGtpLJODCxgKIZCQ9hvOelaeFSr/GoEW93eMGKqqdbjxAAezLvsSkUAY8
FG1W7AVco2GmSSjmeRcHwQgvWyfRgnohqRFXYFzuxX0sYRxR600raBRGhI1E27Fc4Z205oqIbAJQ
tbuR/ivc7lRTYdj9H2AvTKjzysrcRzjn/YCab/uz60BQfbBbaHrMnfN8ain7aZY1gt3CPmeBIg6c
fORGJZCkfVkldCO8oEOGskBpsoNrpju+549ZHopuqjq9njEcpiIa7es0CGI9s1+FGrm8bMueiUGl
IRf7CtNI/oHczEtG3tiSlSbt5OO8kGQXsXF5jvyS5QVbyOqaMwFpUQelydpRnVWKyQLznq1knP9W
gzoNCAqiTT7t5E7g6iudHqTP6NXhRDSa5t64lVoBDyv4SLWTr5heAS183ev4+CZyxVq2P2/ksTgX
MMSaIJBfYkrhuXsfzgOHKUMZTbw31it6aAzHp7HK7P1Db/lqojHuvz6AXaJk3yp8+QU0+ue9EbFN
gVoBjNai+VoRtu5QrTsYWSnn/hJm1MwFNqjFyeV8jZL2L6awpZ1FEAfDxg8Kknmg1H9tD9YSJQoL
DnPio46g0bs+hNF5y33agTwZDvyk0XyMcWjf3CM4CtRLkbdNlt8G7t9n9P3aTQVlI5uyk7Eib8Oa
4T3YL3ar4oPzkgZ5nPcrJouRGzlxY/5NVBmp8F3OIeJig4acrbsLgBVRvMhhknIYHMhrFhBj5GCs
cJYJElDR5pS/6cAgIJEITxTVBXAnaBF2mb9lrCmqNh6/xai03GrqcAapXQSisSy1fahxB0Qo75UJ
tOWvlTGvpZTQYS9b88ez8balIlYHGLKDB2HfIO5+Xve53mD+EaE2MN8AS0+C+i7aymO39YgO0Fs/
ud4O/BZ0K3DBLkJvZuxNlIBWtoGRskJ8siCvUXlNiTRrfxhbLNeZqbSfyRcixRFLKm8G45lRrxjy
pK+6yL4xU8JBaHscnaPIQAvQCZQ3hMDLzc8B42lG4EAjot2xIK8pOKYOqBcQHM/G5kbfwGtcDc80
7AF9q/PBqT3mRn9+oB4sr66DulSVMzMJu3FF7dAeOKgczzQ8YI311zTvIEUxXfWmEXsxqazYsTNf
iLSvep9CJ8Nps5orzakDw3Z4A1lh4fIu52nR+Uw2vruw02BMTCk+q4FtE9WUuuwmoOvun9/JcjHz
e3Ws7djsSGGO0t7T+BnmOFyWqZpaxkMhZoROC4/TnfRSOSZKQx+cgRjrzlMBdkS59DrvdW8NA87z
kK1IpkWmBnj7SlJnX00vzA+iYq1Ro6EFA1xzrXqbM/9Ib0f30+WQOv3XnfsOsDz/BLP2o1D5U/p0
N7/UJ/RYG6IBHABIWf0ow4uB/4sZl9rBkXKx5DRlJXgrC4qRK2TziyM8Ggzy4+HgyT7zZnY7aakx
M2Wws2Q44B72+En906ioYkPqIE0IwHOXCwk0ci9c/oTXJzDnwe5mrB9YcqRlE16eo1Jj2U0ANeQo
2jAOFyEDgZ2aVlN+MLUJ3C5f0dCwbZf2VA5QqIflCkyU2yGiy/l+rHrXtv8CeG8R3Plcg6ZEdAcj
D2Af7/IdGqVuMR4JlV4MzAx/cVTHR+iECTFTewpuHvmvUPPCDSfKMRJax+qjgiym21q7+CQ0Mo68
MspzQwwC1cmNvGPz6fgZnHnNgX7mOHoCF5IeyFrbc6YoqVXTJxRR05EsPMYa39JeZsw0HhcLXSHD
o9KhKcKw7Lw9RJsl72FcjJ1te8fczIdHUljAGgGFkH+MZwQCGX65A/lZ58s6E2lfhDGepSCLVUtc
4naz02vZEiWFnu+J+QJULEzMvtwvkmUyq+kdnWE8kgPWZ/jdH8ETOO2E/+vXd+yUW9FgS5oWhdl/
H7KNgC5w1euzPOeEyEY2GSJHsXGYMhhWoLo/iwIOJzKiHcbCwQ0j3sWCNaVDV+l9NU4a7xWbV0ro
ouGNTF/pfQIP8IDkxZrq/A/aFNjf1wpTB156cytF/JbpeNqfG/MwhbxrBgZLKktIkoZHe2vsJQXX
FHjiDwtcKPVKn5i1hiDqkk5YrJnp1KGMNY7GhhD157o1jB56ip/GdatLSC2a7+s+Yy8lSQ7LTzJX
MbfFk9ylkNjCrR33cep2/e84fyUe5bSM42nGOUBNE7asnq5pvy46k9lft4FXHNQ7He1WUNgCu+d/
3rwwKRQOTVyG1xiuGY7OOvYXFQOk37ntpqOAhUG4lBWIOgonWOmFanKbUVOmwpCdhj5Bi+0FEf82
wnEKX4hosfz8gS4CljMZ7+OVHqrMauDNJGTgMVDCNOS+tXJ5yBwx/5fNGqE6NhRNlV3toXUyDO8w
XbKZ8V41OTDK9U/SBIV/ljBecZerpuz9gc9TgNrsIkkQSkH0s0Xd+q/uuUqdq7ax/wMQZkUg2pnZ
C9sNE2SsQm6IzDS92yQiqbPPWL3SpCT+TPxbrsY5fZzP3pk3rji3y2Qu3KzC7wC6Z9lv2bAmwsEE
PSdDSGF2v1o7zXIHTFMfXkSO1YHzy00ZfbJY9vWtyjfaGbWnDQv63qTHueBni6rDLxpaI0VOTEtG
moCmrXL1FTxBTRCrbfNmrM9rwzxm2UsDqYkhQjJRF4UIkAtzNhuxpgqeqeHRsczw+6gfnmXP4+2e
GpxAApyhsSKQT5QKXJeYsIGZRsOPnwdEUdrBuiaPX1sKKC+0WDuaefxxtZWv2ceJ0RvTmTIzWMC5
M/8g5dAvy35NKznWxCnpAGJZrNf/KjusBCwDcOxZUMuw8f8xOVYyPfgX4PZKumE/VBEp67WwjkXa
4mnqMAbA3N8ScY5xSU92fPRhiwe6xrzynl/upnM+BBsPfTBlDDRD7wDh0gYsOWVOpSh8wFqsxypk
PgpJJBsr9Ntcw/c/Ycpm6qVkyH+sRrmM4nMRQNEg0TUI6QvP+QKzQyZyD+VBHoheBbAqtUEpfFEm
VKS1Pd7qB+EWE8sUEMk8WKyi4NLEnw76TBcCg+Mez+YnUw5hGWwi+1sle9u6d4Jp9s2UbVhoD3XJ
HxvMagyJBhpeMK8WGaG4pzz7K9uYlrQL0mZK4NTNrEB6VnWyjZ90P5Nn03SOcdoJvG/4oQ8NRFXb
W8cOgCREhvOkMNfYfHod84ukfK5bS9F5ezBwZykczOIIoApEovfC2uxTjSaCztm9qziYRPpG3V/n
EsBuSU3TE3Twixq+/Yy3IVlj5jvcqkEBCqD6tf/HFrD5GiZ0KCrXCoVIiGRt7WPEuc1RsEtcEcAS
v185HW0oca43NcyX78mrlq6x3uRFD6J/cbnypR4H6XCJsoIF08ND0ZKwCk/AU65eE5aGuOWSDms3
sPyX5tl8t0rKrCo/sBCxaIJ/iHn4EexWSUJ2OdNNFqa8YHOehMZelGLKb6tSABnmD/4zysCm1PDD
6DVRZQ6+yLvdyDLKIyj7nwMC/oOO2cLTvBrNpiRp+0Nj7iMta79uuQhdQ5cOi5jaJ2r5peJ7sQ5G
+ZSvtBBi/jJd3Mjng0kjhmFi8xZD3/PH8vX5qFnXdrZpoYojHqb1oCjHTU7xYu5bHJoxv1fvTUU3
SCx7KNJ814c06HAPoAybDpxpadPuWxTBuimAenWEgUNNzLkMlW0B/ahMh9ly4TnwW9zycFl0G0/X
1/2sgpc8kbPsg/wyAs9szWu3+o2jiOuY1O10r9h8qKoS3gTpBtuc5Wh5Bw/z2CPIj8PXk+MZ1NKx
uVq4B86W1xetF2A7ay8EUI3iNDkg8qE/N6lJX9b/M58HwXoZDChr2Ly72gfbiQi7Ryct+Wbea3C+
Fd5q1m6RCFwhxhIfZRGmxqU1eYlnQS1tMdwLr1zlxN9A4gjNaOyfveKzqbNb6hFCV1fjCRobX/TK
4uWjgiBYHhcu5IflcHjZ/zh+B7EfJYRJTtZEPVj3RB+C+RUD+n8rBm6WCyEQeJr/htUnxrdrXDU4
mkBSBiZkhgqtKS4b6ql+p3u4uHmFFuJcoiEinUjawBpuU0u9wybSnOuob5uN/QSvAk1giBN8KWLI
OHQa2vy4KnZ0+GwEJIwsudoHrwpaaR98a5CahbxYZLa1mZ8xQHpvJ6w5pTdzUeSSdicELICpAGWz
6aCpATRKko58Rz2hwDBBS3UI7Kx1rW7E+d+4EzZgULymSSPf0N9Kao00067a4Ycn/tbJmx73Cl+5
qrBUts2tR8hKLUZbzqx9uOtDpWFNqc9zWz8CW4zouz9QOsc42XuzCqzuhJO0AQzyoFsz7VCEsmlv
7lV0Ufh9m2Iiw3YPDGb5JhwQ22qQdIm118OonynRZaO1GYW8Uo0NdQ0ghwWgs+lxHceXlUaV8Ta4
7VTJztVvHBR7F5WpBvTmrtjFr7zqjuXRP3dUjClt1L6H6YGv7payVVr++UjcaUJahHSlKxxdqDZQ
ObOv7mj8iNE+APtc9q6FwOSkWVNqTQYbwa+Scx1Mtd6ix7kqPZqw6y1bdSJ6E32cnfKOPet8/V+z
zhty9PH7IDbJVMRMfnVjvDENOQOVrCVT55c8e6jmgErmYbLh+gSdWWS9eQo/usMGCTP+lK6SW4JV
4y+I4tcFJ9fj8OfNN7wD8nDzwQn3bKfhtqUSlHdosn51D3i19Di02c5ksxLeaXRmfzYlHS8fPa6/
2h2aDkIvGQUtQ5TwzjSrSVNnzu28X033eNipTWgMe/+nA0uzwJ315w7gQ0gsKU9kcdMqSF8tJxxb
oup+dLmlJB9Orr/HUauPzju5uNq9CfP/lMkfnG8C0MxWuJYK1DEbkQl1w33YoPlsXuc/kb06zgvn
6LADHGBr8u6xqIPbuumKDBXyZrEkxNoGX3SdsHER+N/0BovO59y6mTCDrr02OHv6ZAgZMKf+dLlF
/l673gb0EthmXBwuI4FUN5l3ssv2C53oKSga9EnsHjnceXdJBfgo//U5hoKjlmuvtFKfS9nBpC+m
V3ehel9ghd8Q+aL165qZ5xOytn4rfm2NwS4HEyuCBKYWcCN8kxsszlEDpWXjwyym/mb/wK7Te/CC
T0oAGxn9vMT7k6Dn2ApaE5Phw5I+OwnMCSxnWaVxoZ2h/BVp8nRG+IRO+YUOFPacuLX1O6KW+qUs
DvY9AVAtiQ64NPG0GOY625pip3XTpgodtAASkC7xXZ+wyiXAtWa54hFn+m2PpkgPorB9xHaoMKpQ
pTo0rl2klVSip8JN72YXir1lmYNrqYlg7rKvA0tXWCwpPaESpw3U0VwNEPDVVAmtBrWUDdmwk6LB
xJnpxrEzX5bQ/tQf7bGZ8soEia+HyMlwf5MjZkY4zn4NgYhmGr2XVJ3EwizaDxhUxnyYKwrOgQxc
9NqSYuJ5bT4yh640bo1NK/aKT6PDtyfEHGeGBmK0uzKG+85PtKx4DV9qF+xUiCqEzK5zbzGZ8d4D
0td6QULokltW7wa4UQTK5n1XEuIOnxCiqyRORstPJ2eyUGrBqz0PxZ2lNahR5YBWwmM2rLiUgj03
46Mfy9Y/KYjqWAOBFJAZvJMLHhl+BjdBCoD4XWoeAts72N6MKhWFN4/EHkK4AXgi8VSp1AZX7Uog
DlT1gNJnTCP8qhj/Pr/2XqSmnS27QwoMN7F2K9Z/zC47Rv6rI0eWIJPgwOzD9K8iWuYesPRYeta5
nmo7MbGxw+8S5/wVXiInIP4zqUBJCKyh2vmuOVXU42QtAZ8KKWZAjaVR2mWFbZJIROHMTAUiFKxV
HVNFXKjEXxz9i14UrOz4eJ+yF7Lhs3Ghfwl1V5Q+RV64mAaBqb6lSEJejIlnkOR0rgAzb0/k/LlO
9KvEPLjuMjgpgW5ib3xgmcrXpVg2mTMO7YJU3zEE+2atbAF4ukxeiGHUGDtBAz/pl3ALaySqbs9w
BmVlFgrgTHyY/fRPVjpqtiPPBcqgpcC6hI7JoSGH/xCGutBEAJNpinF3jtMwyL/1Ug0CIm3bZrql
J3NnQ0VIt/L7wCLVoE2wrMg2DN0dmTpiXsKC+51lWLGSPL5josHUAwYQ1LVTVxn0Yzw+A6s63JCr
p3ZBuKKsYEzCCBGgSvs5sT9Imrrk7YTzosdVHwlAdlatCqAtiEmbZZJn+JH11RDElgF8RQtOOCth
qLrbobXJI0qA8t+347oWWwFvQ/tXUDffNwju9Uqu9XxBz7kRXTvEOb2qMs9D9L+pdRMFj+T5J3c3
bgodx1ynW83d+4+nA5a0XJRBxXI3jIiXqmd9TMYiRhkLufimM8S+g9w46Hlde8WwM9dkS6bwEKs4
ByZW9Z7dkcfxPm/9MLqqSwc6UrhzAxsubJD7NICSOTlWmj2y43Rs56FECqT79nO8ci0iET6jmsoJ
tLHxm+WrT7UIaXPBcSNdOGOGYuUt3yHIlUJnnti9LR4qUHIwQDIW61fSBHKi7BvtkGEvPzye3DfF
1mhMBz65onDj+DEVhmQoi8YB7lgv2UXA2SAH0yZNrBOhZc5hrsSoXmV0BKEd9qfn6aUyBNFJGSqM
++3Xz0LcuxFophbu7qrPMdNaCIW6Hfz5qhfDzdnCdknsZ5/HGMUSX17p0hSnz2drFIZB3T0IoyXq
amD0FS8SHfSL0xsSPUXZ3TGCiC8LOjDi10COObUoi6rFBGUC4gkywwqzguFhH+hFjN1tjThEZxV/
ZpEZcFTUizK9oWR9DC7ew7I5i8VI8YIKmc8D5IrI85KJB1MV2QMhNsBAf/Fc6aYBobh8wEspnbOH
K8eOcRjhWldqiQz2QSe3qN0KNzTDjhwq+uwldA1vEGmeoPlCI9rsnyI60JIdMJIA6ypWv88EBhW2
XscWqXdwUhT/K6E/lgUZkOWsljf00e6RTYWbCYg4FaSrQliIADCHMJTFZEmrvsMlJviUoN4JCbLn
7MAVHGY2t7jMFNXx7MvDRgRqyoAlFaezPyyMNC+zVlTasGikZJkWok45dXD0LJcbN0xtmlY98jBp
2c708MD54r3e3nG0ZW5HwIh2EXjuIMbDWKKWC5XpBDQyAPQ68m7uGkaLhlPTez3zXIP9pPPk6R6R
fApv3LBs1TgCzaJZZt9CPlx7uWZwoBBh7SOAFcIvjAXwTk2egyi/LDi7QuLC1yxelyCJKdNRXbXq
6lVw+DfHUMNpq8T8dV7ge7gMXTUDSU65oZSxI0OkI5CzkQouzc5sbHBL4+9TwYE7ifLzGNwPLii3
CrMFgaXdZeN6DgB3EH95u60rFNECQ/BMopoz1Ev1j3vYVBvgxdJDilX9HN26ULudjksiIYMKSS8R
boEd/h8uKrrRtfl/sIySOKj9odPXtAC+R83Mkn/4KmhGQJBLELz855Joy2l9kOvudttPnMlon4Ys
ClXD/zfk+kJ1R24EO/iI6JllngxJp76q7OTaMdwcUwO6btD/NYFfsHSg6WBqQC64VZBbZcNmfccr
TpHdUkKmbuRRJ6onvcFAEJ9oGltV8CQ1QUNeZZBDyZxapgapEAi0yu/QI9b2EuFNT20C19Kgypyj
paFvDNoqKtHVnZqeT8gRoGXtTt1WPrn9gRHF3pZCHGBBRyo/1FIutIDXWp4j+V8z8ljbIb2mAcwI
2yZRVAFHd7amy8Ny6nQZRuOD7lQkOhd8vgsFzvQa6/1QpUyPapUFyeOesFl1agYolgs80MtXW8dz
aXvQNAGm7Rd+A+6Q3PjO+8sPHx9P7o4q9MHQfBLGLggCdrkNcJ/8vhV4eS7VObzGwXLqxS9u40pT
iA/WvMmMY4JmpsjcuuxV7jQluF12EB51rcd/9nJ4mzJkbOO22bDvuuj6MS7M3RBbAmsSjo9UeOBo
WVaPrE06YKHA2Pw20rQxsDrqjOYzRK/JLzrlFnPImulyYmPz251w5WTwXCatfjjW9ULsDe93dD+d
R10ykKv7qg61pcU6PeDUCGW5TZLvWgpufUXVQLqsGWnqam8793Yvii8IomkXFHAqz8k1KWoT5H5I
ZFthJ4Nx53OjonBL899UD0zpkwUC9bAwifn0c6xuA65uNM/kd0OlxcmhxHjLJrVzGEFmx0+T56Sl
nmEZxIwaJdtQtikcDDxhelMkXlKfvCs9RT8m1UQbNjnHIOQf5lfz0xyVnsqHbJx0FcA6Piej3Yz+
c0qXUZH6r2W94SGnqKS4x16UVFSsU2dvR+LN2991m5kcH7ZvI/48H62ZTakTRiogvJ8jK8J53bNb
PYU5Vfv5mBuSKOMeT57V7p1cvuZzn5t+xpUlAn4V2ksc+GglivWHUd0ZrqajiNHShadsCdJFzEzg
7ALxbmyHphwfTPPb6MSCCDUR060qrCvqOAdtVJOD3hzue3QjAfcwsAyere9Uew/YRJwZ47t1yRO3
y6jPKzSGmLnjC/rYM1lNL3DNoRLNwwq2i2bnpYUbmCmGXcY0WC/HsxLd+mevmmDcMOseMyxxAqSz
czxs2tv1ZcdX+kIzZZh0RBV+FDxOrQXt+fRJIHoYVDq3sW/sRmorq9sAWZtI6qMtQgIkhguXN148
xFuMTWzqAhIQxTd2DI0uSFUiQN11WD3gCzsPIdX+EJaBIwd4jlN4Byo8dudOMuuomJ+ohGAbBiKh
g9ia4n3xu4SiaJDm/B1WdpKAx8YB2NMIKf2mZkAmfhGY5GWIBoq+14vtnQTpnkDxds4/Kh6sybvD
ebNpcKBaX4xuYdxNe37wylHQijMbKw5SOPmSyGVU9byynatN2XdxVQyZCt5JjupuSWJ2acECfY4C
QzMK4J3mxgtJJR1A9SmSWYqtUv1XQpsv/W1aY2FbW2RyH6sbQN9MMiZp17BbBFEIHzlsIUj7ReGI
kaUkNGz70nRKGZbSn1p7f0f9o5JxlSRHLcULmGL/O2t4gZoj2upykgdrywR0+CTdykyNJf+NcEg1
vXVoGv40NrSlCYV3Z3TNx+FW/sdDRTPh+WH4dqiuHhDpZBgKe5V4sBnjcOZMR83JmIK314IDW7Cu
wp2GdJ2DmNO+XnSwKUVz0hhBQR6pwYtfKT5ud5X9O5FzUUmPbPQv0Gh3ETbfzUiRzsxlnjLoB1Yb
4jtEDOfiWVooQl/Dfu7mpIyGBx7HiDaArYm8vukbN6nBFBlHfrpBExVGqb9a92dwVXgqo7UWSF51
lEFD+OZCg9uD7FDhMqrU52uzAULNwPitq6u/O0z5x6eIArpO10TeFBJlEtS8883SF+D6P2OHHP6V
2l7drN7pa/KTepIXzmAHQaEayaZdKfCIFayPpGUmpx6qaWCQ4YGOIWoFRY+Ubznzledd/nNn8Ujj
5dL2C9Hay9n48o2XlV19RhzXpNOYOk272ZOFl/JXZm+Gg1bZXTgayuvRdriYtiiJxYSdMjutVoKY
4k1yFtQ+ZHuzB9i3yTGNk2856TlmgJgA5iwyyp4CdclTSIeJRKmcZqwhGWq5LAo/ARtdmQxqknQ/
Amtzidu1xrWg2AobBKABCG++8PRPKa/K65/qDtlQC740/kIdoh+jpvHcQqHqKBpNwBsg7IT0Kw2j
vHgL5ysoGlGESObWwtzksOiVnYmcKrKw/+dlB9WVbr6gSJTzjpwmutZj5LzU37xYu1dMYOxYaYJr
+8euL2FmMA5nUhCkNR02NbXXZGWXqisJ+qCGGDLJKTP1yw/jJs96MzbBq4rsVZfbn9CcgMz8C+aJ
qFntgt+euap5xalF88xP5F3ak0YRXPCwOnTQynYS0tB/iMsEpZpdsqrMsdpwIlHFsbxDHOeDcsy1
Fy8K6JKdGrMWVU4Exe/KzIe3Sf8iRbF8oRQecVTG5Jf4F9RxmcrHHCToZvrPpqWLTaBgX/s7x4/9
4iPsof9na5894xbHWjAz1p/a02Duh3GEgoB4kHu+ri1U0L7K4MzesHjJKELCKCwd4OpaJ1g852Aj
l5Q9nIXATH51i8+zHqaR1h+/wl0deIiBB0HTqztQbv1nJATQgPrRgDiSkCRsxrbVzWGru/cGFZaL
A0aeRLErf0gW1OE1d89i32uokiTPK5/t330sB+cXnZw8Cov1jA+25kRMgVtlHJdf2kreExXL/oK1
uoA/naRXlWa8z1mh4Asa5pJDAMo0qAvpYCXOGyzIAm1dw22YCXpXxKbX33KFO68C6DYt/7GRphhG
9425VE5t2CsVMoWdCyAISxqqYtyv7SPnYmQM+n1oiKQxPhG+yHkYPmDyWP8UsVn/5N9sKMuUt/89
EjaXhc1r3N/oH8BBssuNI45Fwnh0WL98x017Xxy0PFrgNNnHqNfOYuLYkzq0HI4HVNOxOZZzLyf6
lrMonKz6qQej6PGDAwpZdq6/2MtjmlQA6xktlzhtfAcsfzWqzeciW0KfPxAs2PK0TkdpdAmnjf1g
PpPG2Xc/uordqkoqMEiTy9BSRxb/VsjlXx9+YSr1OqogyuoPl8mPUGUCCJx+7wr/hF3WammNNnwG
JBEzogPA2vUlAl3uhP3ybq5JPpSjsstJ8xeMQZ01K/FIDIXQPhE4EXKVP2spMdJEvPvSp5cIEOan
gPEVh4uMbEQYRxOLrHZcC+vb301CTxREksF9jIny628ZyP3G7BNGwg/E68W9jMZFmi2gq8Prv9uY
c3Wnv+d6RvjZJsDat0hbYfOPj1hj9f16+1lEp3IHrw65+JyryS/qAlYKCztiNkAtCUHW6TSuPXrH
tDizulz/H+CfwZdQxUV/m8dl3Y977+F9zNEx4g1XrLSt1Xwnktq7leps09ox/wKqCYZZhzmBplxn
tdJusZwGhqaSFOgFDs2QFoE934fc0RveJEdEz+HWmnUgCoF0+t8bBe7HzC8zVYpUn5bHmNg2i+2o
Gw1RBZmXoJz1JjP+kNakKvmqbQ6VpZIYbMsVY3CN17SDY6smYI3Lv41HfeHS3CcE1q16IFI8zHKt
9+RhVfh+H+z28RpHMJfV5ygBGXYaleRz6YraLC/qTa5aXlnLkxUfHnam1FX5GUProTXO0+2l+QkO
LBLsDhoXtC9sQ/mvs96ehuImij1h8gvaGgyL9ddhJ4NVsMPJFWncYQyuolRlGuPZ+KK5dvT8R6SA
yn6xlrSvB4lhtjfmDWV0ACj+c9Q+sWhm0dVVbXGIVDxZDPeMpyazNTc5+fSnUenp1oM9cWf+nVLv
/TZAdvIo3KlSar+e/NzM0sau7d8EgBVU8ss8av2V5ghqFV2VUUj9tYJLwr2Yd3UAxVaz194zVa7z
3e0v1jAR22gtVDadc7p4lZiAS+HckPe/W1/2itbOQUrmZtyr4nkGAhLPFilxCcT9ynSw9wfBRWbn
2v5CLzq1A8H8u6hUb4J4En/q9AkY28dodjMPzGOPcT1bgFNU9sMdrzKU4tqn0Vi1epXI+r3giZGY
47h8IXuAkfS71U3yT6aGJg5lXhtkal5R/dit00H82RyoPeAToCd/Tm0ZX6De0jp6o702Y6QbSZlC
eK+8VyPl2KpeeFEYhKcgDoUSkL3cd/v6XHxA8xj1tWRHXltbJTu+KtqTs2k6MaHEVPjodaW4bdzm
W0gFFNRD2eXrwoTi/ltU5ZI8JgpoC1qc/qGnDUqBXNAVLSZE9M/sLQdSjzn7b9CMGikZZLfhopK9
PTetGXf08lx4QCgSynKb61VwdtXOoMusvANVWgL0Nvu6ZqM2rTbQaT0vxh9NM9CUCg9Ooeliu6hH
s7smYdM/gy7An3MIZmxUzxHODrWxOJML4myi88m9iCRVm0CA+P142CoCUDT0/BYIBOm3x5cnkoIz
w0xKCO3kY/Hthxr78lqXTzwAkDzKEK6njAVZPy5MMjUaWgJw/jt1XSTY8L/D4rktYZXBSfFkaVFX
mFJt0/vN5WcVHW/44HhnuqP/dELQ7zb8mLAHzW4bl4r2v4dN7Qe1ujljN3GuI3nHSPmEsjY/eNuK
G8ao6BZn8l1syG37AT/VnH7isSyhF0FFssqlMSOpRV9yPph36cKxKl2Ew65maucDyjHh1vX7Ojel
Lz8nuPfcRAD5vWHhW6P/d0SvSiEIJsi9MU67MC8kGxMv8jGAfqkieK5DyZO2iNl1GBMMHzy6Bro9
i+Z/ppxQiF6FAHUB/neFtzTvdsXF938hmJtAXm056F/O7nNv75AeAoiByhP0cxO7ghluLNRYDdKK
58BAf7/CuimmhHaoPW/1FS3WxcFfhhl3eZtW8AydhmNlTIcim9U8eq+/MUaV3qocr8PtyO4ygoX4
k35iB66TGA+rGU88F2m79og0fm0wMoS+q1kHHFF9OPYtczH68eft8aV0wZ2kNj+gk3BooM99jORc
8Z73hrEzr7seKLV6hXlKQemaXUEHM6V2bIz8w7rmqNbG8oSrpWQwDQ8HS1VlJcLvFC4yVGH5QaTB
z3PIqKepLz5hBucdRAbngUlTyO2hHgg8itdrM+z4oiqRzSDUVZG8kx6wcsmxS7q9TPI1MuHxD549
UCL2zDGb1C4sME95G9/WHyDxnUI5LtwFSaDh5BqQHXuYk4Wai7JGTatbGFm4wGUXFT/4FHwxAY9n
avdT6c6/tLBO0rL6F20UycBbSb3TTWCkVmqSmDE68v8CozWU11yCwl3mEZFX2fTg4EFBOaG8nwZf
QZgCzVWmqlSWq3gdjqyAHv80BWS9TMt/n4nlxjNDJ+rtqYQ7ShIlSTjRSDTYl6Qzlkkns+oGDy61
eMegnsz+NS6fB0F0SPXQw4sachgumtLpwqYiR490HPzikBSS8drhfhwF0ceD+c7V1+UMKkSWtU/7
/PUL/VP+07CvBdLnf+0GrIY7lCUPqyvl2Z4oh6nVwVb6Zp8kMzrqmO0+DPToXRJSuOLh+hh4VMk5
rs+c+4rFFs8RQeWXQzLc0MEHUVvdGlD0muJvrcRU/P5Gu1iSWgT2ZN13d/9LR5kFExHAzfEiPU9+
eGNvfohpKiUTOzWgLIzGyJ4BI61kEURg0+2o07cuiWK14JzA/FneDIqNtUncFaHJfdAA/xyvg1hX
b4+fF/vZ0jxshiIJABChy1APftL+M09HnoXijEWSUVbB9EX/kOmz1QW8ARVdqDz0XOhlwokhsIDK
wJakW2+oRaffG3XEGWCFffJIwby2PCTAe0VYi389ksGYUSfLqyM1EMsbPUidVUl91NqClBuUB3zp
xgNJlXnfDpU+L7BN4BTexfjfo+sOvQJRx9iXtkSHsYjZZGb7JOw/WdcPJ04eQu7EyhGl2BepqQPh
l5LUXLlbkhg41iyQq8KOoI3q+yxsCW91tAOluKbJI982NpJjU8SKe14jQJKFLJ/kXI0NWb3L+3vL
O04tEtmPDo9E5xaF/zRI34qY2kZxupyQUt6B8rWxZhFt0VONTsNrxiGeEIUducbwTmom5rJLdSul
vewE8ISSY6v+l2dRrWeKG/NZPGBDRLjd3+4gwHsYiDttYJWpJeK4ItWcUYe8IgcRNFm+x3VprS/M
bGvDJwbsK/BBRKpfPXIk/AM+o3ra1muFw1Tg20utwfDBb8IWPfbwH7ARd5OEu4Wm9tRDUoNOleae
0Snr4gt2XitDihLfANh/mMIxrXAR8gRgXLLBzXM7cq61dMdaaeukKQ4fFdS2slNdU8HfrTNtZ1E0
7oLMGieIfJFWQe24rxvJBzFsninim24Renze5jD3fK/BtYsCsJPkb4zsPIq/DGApG2oPsHXp2PZg
KCqrcrlMq4VGemdNhC7ZkCEZjxne8VouUK4FfL7LhD1JZiRnndhso488QX+xw0CG2f+XApiUHRNp
EO6IqzsnYKgydwTIod6GHnP70Xm0Vs1wg8+9Ub1pFRq4c/bhL7W3ZrEVE+6iteI8Zv7Nz5qtbUmh
8f3SeuwkHGoJzhXPSkKSebPJAgSAPDmT88ilbTg4Wu02JNP6YDKKyVTaaBgu/A8oPSHyJDHljlGC
VfV9q8y7CUYE8Qvhuth99AiQQo0kVbwSEqDf9Jd0nAm+2QYlK8G/1hRawpmgSYxQQQlXDc9TG7Po
6namdsq+lC3Yq2uInML2Gw4OUp6Xml/fjwxgoY6CP4M1Juy3RlGlCrGM5LliKdE0msICGaXEFC0m
FdQ0UFgOApYivBt3lFJhouXW19OsiARtwnDzcfh/5EQNrOJBPAE8D146jatTy0OGqpOw6lizYWKS
wkao8RshPAqY8SXWLwPnBgfFAxCEO9qHn/IEGQj3bHS+AI/l3idyV+fxxorhASraES7F/tnC025K
4jB0NQNWiVXeIW2ZsYfIitCE6CkFrxW3Q4xYgfHJp82pL92ykPt7Ev0ZoGfbCgF770m0cPRQyhXb
fyQmQlcRMQIe5hkGj/i9788zoexDKXyJGgn7uEYMQbaxiJ2hwRKCZIajL2rPHoT9A2okXMcUTKI4
8L7eL0CbGDkZ/6acXYoXnxoHK2fhue/NzfSVarr732WlU5FUKUsJ+31HxPoEiF3VOfbL1uhj3I/+
Hxlz+MsjEmfRe6gMx+o0A1cvDJpk1Gvn5+QbFhZJAgjJFbH+b+S+UPNaSZUpQodA8qJhrSzbbw+m
sbuxPFj7R56UOBjWdj8qtti8by1Ihioh0Fvdxp+zJ0/SL3UFjNqXmI7tdR9/V938z5cAtVWMo8Xo
wO8zVdydftqBXf3+2hE9E2GWjlzFWzmFEW4jhkkGGp1XD7yEWdHgjoy81MLavfdWJYwgoVZVHohi
+rNJqCjb13He4PaD/TXGvbpMkAVqiPN8pZfhum+mnHo447bOJnRahWeH3FjYNuy6DRUFF4nbdd8H
zHuC9na6lAoWK/a9vFsfNqGcXuIcDDipqZenJK+BChF1uJ62Dgv9qv63KFmLOecgQXhNXOMOgg5Y
shOkMuXI9a9hZWYP1ol57LH4XAz2LPaUevsD9j3OvXgaD0HLgvntKQULa9ZTk2oBQprD7kMP44RZ
4gLGoLWmsvWGSSpC7LfLkEtFSVrOPBQqhoQN355MTOtPff4MzglOKWLKfLeaPVM54cB16/ZtFfgX
HkxUxuxuM6S6jM2tY7kfRoU8bVO8Rr1EAzKThxK8TocJBkfOQvN9nzWzMnG9KbiVCwZcubFDxlS4
JUtT8NFCKOyz1ZIy2qPDYt26MRlEHlq0wrKVdda2GmX1uINEOGbtnlotYPCRYw/y2hYh0sAFfpPm
/sic3Ucfqdr22X2w7IjHd+69e7qfFv94q6pMUvF32+kchFlJlittDauDQWUBHg1YwggmoI8n7hL6
2nqywQgbPogCGcfIdsSZZxHjT/xzSDry3RXXKPCUh6t+5un7dbN3EndkY/Spckv1YUVOVS8U7MCB
7eBH7w7tHNVb/utTcp0iEQwWUPXBk+aFc3q1MBHwhostUqBBck9VlnWPJjfWzjXa3kxvlisWEBHQ
QQNppb95c0j+qiVpL9MQnFsodSD+4483GM7Q0bLHahooUBUTEfHml7gGNKLK4taxZ1/OyOWso4Tt
+8mY7zp3xIBl24sXmKpZ/aKDTZnuOj4oFZiCT+bdKr3SRKTAWnZjwgUf7hQ9RYwjhLFIDTFnBxr0
vCwP1aC56sdrdXij8o58n+Uaa81IVTJzsmxezGNYDn7NBbyAcnQhzSVywVpTuN4YB5mBgTDUAdDN
7+w0XYOxtmIX1016buj9nnPkr/uDsozLiZUoF0el1B4mof22d0H9F9JJp9oE7lqcd4NOmYT/Hkpt
qD0xLDGyLYCGyTUVuCYR3Y36/OZBx++bHhgaP5tRumxm3id7UXP4EVTAF9RdVqoMGcAgdl8dT6tu
+b1n73LEWO33VQrZDIaWpAi4jbW7r+JGdcE6j81oB6L+RxdXuP31Hv7SCeyKCLR4cFNt2hnPR1Rc
L2SWmTKIRbzd2C3uXtDpsZvJTzheUQPlGLr2Akk2ave33blRWLvivEaDMhO22SlBrBEZL9F5k7F/
AEKs9zm9ekdvLFAZewu0k4JVzD2EtF/6UOJRxeBmOKPa/DlZaA043AANiFlOc8xcKso/11mWTyRL
6KubdyOUy8soCfg4Kl8ZzCmMZZsRczfesh0Qwb8uiNnXvrpdGfqkD51HYbjv4AzpeER2nIiH0sD0
XLVPBocN1knT70iikEANhtRNMCDFw4RfGx+3E/7Zi4tzgeUTxqUaoxePIRpTYZ+F5aLA/JX79pVT
5SfC3LdsWOkm5uuvObugVldH33cmth31r8NzVxlUppCkfm/ixRjMOQI4SZCfg6bJRrhhvoFnfZeY
E3qG0elKGlFHXV69b9J02fGutm12p04p0vgdeL6rYJ+2T9ag4X489bFULVwGtAFrPdZuOPUwp5Eh
bqLYpR4mKjGkIgEyJ6kDiTUYgL6YPS1BFSmgqeTiDg7ERtwpl1ynvdu0gp59sI3xSDxsNvLwF/8h
+1wOcihm2JFC9h1gSEAQvKGAyxH8r8zfvPpeOMQEtKon2pxYHzHUhe6hLIoJkmXypXzkXoXj4dZJ
UTN4PN9iY4+BQDJf7Tdhjsxn5a1ErukAOXmctUw511Lv2l+J0UCgnYSQATmaI609ZnhpIGOmQQCS
hJ6Fxu8Zsg7EKd/ujw+5QcgKnurZl10TibC+MPBceIHsgX9rPRTI0dJi8qlbE6GyxuFNqdvDP9sz
aeUB22zZPKn+ywWsE66++5uAMO12OUGXfOMbpf9fo/Xb7qyiYJM62xkgE7zfZNWBi1PVWTvef83N
O3FX0lAtd+2Q0lZTTCH39517kAZ666bZzn9IoCkjLsO6NJzkC/9QOD2OyiIfrOfB5f2IM4O7GZHw
aODCnGNBwlHqjzj2WOWSYlcnePl1pIVZPOIY0nP/QBlPNi4CGkeEZkq5J5hUcat5HjVs382JVNEC
kZ1YneySA07mlyt7sj4Dwem3BEWFzfe2dJ4v94z6XWCxKDu7kO0lHbGPN1N31WIL1kgCt5VstEAB
841RZOMdFk9Q0LC5gArTv0G4nNlZzlLlQxF/BwHAimYI9an7gZp3WP7HcjsYB6ri92f8D4VVbLod
safb5Ebx0Pm4m0WspIMjb5sT6Q5p7kCB4VtnHXpwFfPHVq0M27pKr/n0i2GG4s1AEkue+EDfjaBv
sQNF1nUoaTQcpijPKS8v4jSWAEio+17AdoozATs/JcGccml5wGUlE1590pzGW9Z196rAE577a/Fp
kaMfF1tMQvNG3hpur4D/Uy1Z9GLATLZl2fQRBcS8VDbQkaU83zG2eG15FRY9HSyYH5cZQsjkm+SH
jFil4dLbq9I9HSHSEVQrZvbZ2+ujtIGlvfHk4WnpmjmrdT+tkMoM+yrnoLxVfnVW1iyqaYLYWKf/
QzXuVXSXPrqFf7MYzlX0+hVRKI1oWb9C2SUVYunEiqS5bLezUcqantqyfOZKI0k6gBhY65fxFwQO
bx3kJZ2p+UywZZcbeBK8cKnA6RQnPvwnhlQwL3+7YP9lyeWsJ0pozoS6kF5kM5p1Y8X8rgPAZGDU
7Di+F20Mv9fDT4jX2cJ5PCw1IVGIu3Jw82YP9KOjtroz/L9lIGnePkt/5fuhyEP/KbH9fXT58s/C
W308G8r2o+YEiE38UKc5hmk8qFXv41IuPJQxJBAGghfSOWxLBga6RkuUg7QcCvcggN2crVdMvmdo
bbAmaPRTsjUUBLsXsy6TOEoPiqlX7h+tn0VCBCJwxNwosY1IIibmemw1+MFlPY9Geg+ihXAJ2Yof
MgALIIhPjSBvPFRIjgSmmsAGF31gx5FMh1AVSibnNOhfY4wOrH+CJejQMsARK4vUoPS24UXq/0nL
/xV6iacX36kz/ceTE34EsvkGUcc2CRU5p63FqUoB2Xpbfl3NSCfUeeqE1aYg/ufUQVF5AzB8qsFq
SiNyszIyeuSMpsEHc8C5wNCAlxZBqIL7a1vR41tUCXE9th9Wg3Ha7cl9JKwolAaQh0fYpv3bIGMP
JL6VA7y2gt7AyitmXSSNFvxYFcBfjtSKDDTfkb9RvIzWc58YWEzM0Vfa0WwS0d+14jnrVMIsHpW/
aGTFHPhxoSKu61S+xzhg5Js7uLeNDjmcLowtB6B6V5mjWYTbL/UypKfxFKsx2Eeicr1agfyIVGDR
YDn+mv/VD3/ag5xwoufpdZKrgSFAEF1ejoHvfXmAmW5HchyzYwmnMUsNiGoQwoZTUJsSYe2urifo
PxVqWjoQ/PT3tqLyacDon0QJWzPvk7U++8bcMp4MKwzvIY1qPPTZsyHBWDWo/0SmZWhjacE6Rvga
Z524TXTrU7pmJwWCCHSvHlBgWGnCD5PNvJPpFSVz+fyhPVD6XHF8qcEckIXJHXSoD5LTKbPNHZl5
cj0j2YO/qbLywYHfayIBUy49wbwg10yFacDjrmVcAOxKpIs0wO8MjJdM9Lf9S72K9oJ8ECR7gW5W
E+6q2CF0OR0TgEzoSvAWf3jEgV9nCtBJWuaqYS1OyRUUDk4PWg1DbH8W7838GgenrTGd4kWjpKQp
fjYxZkOpED98CDEUIAGm9Mml7sVDOYdywROqVGYlPSJKFHZCLUdOLuVL4RLRPk/OSZjeHG3KFy5B
+f+aAaTtQWS1SgtBi6FeAPQfscS7B7cg5thXA3rqp78kNPSISw/1BjFXdA9KTwbNsc9lMxIgTirZ
87rN+LZr+1g3pQ3iwR6C3trX7Ne0K1IQ6d4iYbkLKMD0t5HnqLfVMNuTJ5RLPjOdaepOXHc1ae1y
Pfk4eDqtsF7IibO+RXnt4weDPM29N592h1a0Q5d82NbZ00oAhMr1w11BS3K60Km+fzOyxuHNyYDp
0AxWDEkICAorZmZe8Dyw5+EQBqEXUtf2QwZ6IYO1ZMvUPM8bNmDrAsze3Z9J3T9Hj66p/99Qrtl4
LzHATJ0wtwvk9DRNCD1yIitJCzMeIikA8imYoXIWFXqGL9ZYvK5TfWM/x3SPh2qedzsbYc8ssSLQ
przVKDS+hOkQFuGX5InVmYG9gVwC3FXgueryjwDcnuoxhW3nCRL+hHSfOKt7oh2C5wvJgPNiwl4Z
uaS0rHEFPzzmXBaAT7hjGyhVCaSniOwq6R7Ve+Fpkif5I16OijN9GxIj+s3i2/VQIYMyZBAz4e5N
C6pJSoi+EKp/e3rO2dH3gBzRdGQCKxuvucjRL+h9TNYCbwJkFSZGxsUyVzjMVjPlzXXXtaR5iBUR
cY34aV3jPr7u4V2RMG4fzN9h+WylrPdUJ/HxMd3YiXlatymiK9Es1uWcxIqFnTKmYCUgfPM1lu9G
ey+QInHg9rDfQbDTEp+kK3CgLQ2K0ZpbuLffaKj7oM3xzv3Yx6aE2e2o/y2Zd+dsolWJXXaMxJan
B229MBLN6xxatlqAcnqkIv0NqRXd3Ks421fMKR25jJxI/pQ3MudF1EpszJm9/gLCZ0Ml6WjF29KZ
MNm+F/0fna7Gvu+V9UmmxPjXhIJRA/JFaAmHfqkx8fPARsqx9f/mbK3B7v3wOT5t5e10uqEkhgz4
3u+bUlQN2FADJUZbfCUCSL1Kq41g87+NEOmDgZ5DLIVVtxOZDT6OakUhhRx3eQWnlmsGg+HZ+yAp
MuQBF9k/kYJ7EGzGOP55IXviFzMbgLMs1Ytto7F+4kNg+jLJ004J3RoT7YIivf0ROVp1VX2gU71S
KsX5+lhh8OVHAbanwXj1yaZblKkA9wlYKwPvRinB65gtJOREt98LfnDIl8bGd6+dePtyhUnIXdPR
0OuqR4zkBCTXrAsuisFW8ufKI4hd+m+AHV8H9uHQmNnYVTb0+cUSYiK4ebVqiquPVKC05PF8NJRN
OTDSCDRikYfxyZ4e30ZfpYpkXXBUVW80RNH+nYPW3xGTkkFX5JFbA98RdzxUtPQH5iMYO5g1FiCk
lOqOPC0lsrxx8rnXalnoUxfvj95HI3dudqpvAvOlSqIC2fqZm7uhjj+iRuJcqd/vgd40q/OJgw8k
WySbCjQ8BSykznuKLD0uSb0BqKt/RFZRerzFJ+l6RWbgopfM9f1Jyzy3CiAl0ZeNg983fzW6ZOn/
NG6AFEY9sF0rjLEuDTGFTiWwW7rCSGwbs1iYKdsN6wbnoE3QJF6lt90FzjATFbND+SMLStIIWHzY
MWrZxIfpu5vPT2fYf83hACQD1tYAsH5ykKFDOYBB687ZNwT2ur8WNvsGTd+wJSf21OBdjdFdblj0
fN6/A2Owvu1mlaZTafj1UAdQS+Npxuq3dOE/+mP1GHrUKCfR0nch6n25rnLPrbHikunHvwoBMIFW
mqM/rjDntqpD730E0am31rcfiYl6nUYeo1WC0FlZT+XN81AzFp23m8lKRLaXWFB0OGyKG0laulor
H8M8mbWgN3jGj+qxHObzweaxXexn7OEe8BWFntsx14ZJXH6wums3ZFb4blpXGMTZjsbBezmLFq4o
kvgQouqePVH7eCIsJEerwfHrdhGYg4akULwRT7OFdcMcc956lWos42pH6oNA//hhaLVCsW0xXwRQ
zDqDkSTjQjKtb/OtnLda+MM4QDFK9hVcVnSU888TAonUE/oKH3rL15GgYArGyLOfk8B6D/umgCHS
VFIgDdCd3rUrIbQ3XH9K+sKvgUH8vwpvEGkUBvSOAkK7M0D4Bw54yL8mt8WfEw+HeuSz2IPdlYWt
Z++3LWBDKZNI7xqvVQjoUyeL8D3mUuRwqN9BTNeiCyQ6qiTd0PntHyoUNd4sd+jrOZ+bKyxJCcux
gJZW9+Q6WXrBrexQ/iyKaV65MrDtjSkVF05Q5kYdUs0mgE/Qqj2pTy+XddjOaYBufjrcJrpBZFjt
AQcUfTVyF9uE4MKeefdzE0KnLP1Bu3GWUA5gJnWNX2CO4AHQlu9s/0cusGzIcnYaYdH7WNg/JVNx
/GjCxxw1cX47LKb36Y5h2wOEZNtA4YlsWeSaLph2uha/ENCMqfa4i/wxA4TmMloNQ/bBCmyt3du8
q7yCi9qYWotdIodX9nO8MPYMl5HM8bAmS2/94N7K1tJf/4OYPHfeNUvwK4P0Y7PdbV2cxpQIl4zT
/7gogtSbXoH6+HNrec80wC+uMMIiFxaFRdE7WFG1i+8rFV+QQCLcaPfQVAfX1heAdKaCrjmPXcWK
KJq0zgjvzTRfP6tRUOKo4cSR/w+hFAlWNYIN++3SZbov+ZemqLHG07+NCHJh9TgYU2DlS6cSOrjk
WVxwuVjQvyI+y0c+7MJG2/jahApC+CEaB/8kbZmjEf96O6f9TOTEiWUWcZ5nUi8MZ0qrvolIuMPA
bWWPDQcx66RvPx3jdp0oUfZqpt2Q4IwfFRDnZQlIT6zdhOSDXxyxOXGp8UeFYk2j5ajZHD+7Tw+7
GVN+5aWux+dnhsYUfGiTxOzL5NG/HmDi8KPo+eeGAGwI4fewzOU+R0Bxr/jem/EzkQKIxMOjr49/
L9zFJHW1KivWXZwlnPyEiMVkeDW9m32wvXhCqKiT/8Bu5gLnwZaHYg022uY/y6YgpJBDMYjI0esG
9mdZu/T5NZu42qQAWiwlmTaeECXwp0sKkUf8QZo+dY0mvML3qEp2iN5JT79tq1lUZ93DmDGjLIm+
p64O2kqiVV2ixl9Q3rTYag7+/niwSYlpVQyUUN7qMYv6O9wPuMnKtZvxwzLRr9diFr4nWdqBOZAL
6G+R0zC+RmOEGy9+Tkzwpv3Melei+rOpQNpk1CKHdG4L3MYH6X76bVCMXNhwgRCodLJxonO3Cvsf
bT04Vk4oG1JM1tJVuN0pNg+k/+67jhRLbcS0BZA70X7ksso4wybpFGwKDmjbRQlpiQx+kX/6zrxI
9or5b+MSBZgd0uKthHzisNcRbebCiqxhungcN0Ba4gs+nddO8Q23DK7B0VITbAqNmIEK85ksQpJk
Yt+E97tlSM9aCn/E4XsTtnlDLeaMmbMYw1Tnq5b3LISsfuRM9PBE3WgbcNzts85Rzc4z6idcaIM8
ZGaMRNjYz6V9poqZuCqxJLFgbn15piXbV5NzezexNLvKwIULx3ZHwvAR30pxO7xNfViL+wAiyl+Q
ECWAUd8n41zhnBRKll1xfaydgHxBAAcrnP5gYcySeWEy02b+zfMf+ocwnJPbOpzITzEwOQerirdO
7+r7187PQclsBDoVsRKCItgW3LYPXjSoQc2WwKmFNvMS1b8cdeZyqrxSohd/eYek3GccKniMAwSI
L+9MYtb+zhQEMlgtS1GWeA7vY9vpBuFR1N1xi2bcvgu0SHISfuZqBGMUPEDZdFcMipjpWCycivmT
x/Ec4M1rlaU6o6JEf8rpelHMYkl8sEt+Xc6VdBk+ef+Dc/PLJZkJfdfU73Ds6UhLJUwn7I9tKavv
GsYOdcdiWHw12RAKBxc8w6nkg2qOFiJ8md3HkiS7vFg+LoWNm0oK+DPK/QwrjF3DJZ39udSWa2vZ
tn6FNJOdcc8dbRaH/kWmGQihEyVlj4Pg8GEgiSXV6epy9rJ2/LuES0TPEedhuDP4Gh+IfAjWDTIZ
Q7uaAPeZYMWImxwWgiHyL5cDM24uta5+7qNBDhcr1UtOy6bW6KC1/ZKG/XhHlm8+zFJm4UXy/OFd
Xa5am4Cs8Ags9i75CqlDMQtxPpagLKCxwaDw8bgeEzAFHINAcSiozSY2vSn97e/2qSeVX7w2fpdQ
uJgkX19BBZPHFrfDlS7KD3OcBT2hbVgW2UAu79tK5T/5snFMg3aOvvy+ldYZz03ZD6z5T4fduBlX
1YPLCduFNq4uS6F0ugSTmj/HzT8fD62AI0JPnb+DrEfVt2INCGDFdcaW2uT92yXAtf1Wim0GxOtX
DGiWYc8e9i2CeAKQ9eRAaHZmyntXykutLqqUicxAu1rSaXwn7C3Tc7xF5z0CZZYJqVOCZrr5duQZ
3mfdujHLvuKbylS2PdDta8RTuU3BDsuNz2TQJWswzT2MbRr3sd//URn35Ow3oYy5Ueq0OkUssGtK
DxpPyEDtcxTD9dRB2mXqzMh1K9cN8xMFHLX1Kj9IMQQUpTWjly6hmh1VKYyHczq67+ipvOrj4LQ+
Fxa2ftT+qn312Pq8ZKl1L35Ev0RlEb+EtF/eG0y4T+qQPcsUg2W7gDtGBOWb/5dcDEGDq64wpyDD
UOyj85v+R04yQLkjZrfOOt7UT57Y4PnrZHcjXlkIleeQZzC5odOIKskr5fgTK3/P9VeL2XIG4DDf
FezjsKQnHL+76xN3uP0THqJigIpOFBw+Dbo4bL+iStEK0YJanMHhyUlqqFGbfdeHvrVumVcrC4M0
e9Qx879ob7GarBm6WMjHK2M2Hgg4o4f7i9RZ/oZUthYEaRNwX3RN1VSWfkP1kTNhu0N3lon3i1rt
jmzdtLO/sXGkCelCop71p4RhNbutD4ga6Pl1EjVs4WwO4jj/XAbZUWEb4eW8Wp/BD9xaCDRyhWKV
OI8MwA8b7vhwguLh8ae2WCHTK5CZTDXVDOY6EXJCm7KDuQyt9yjynejH1so4rFMbRyN57uKH0qLT
ObnaYF9uz3taN/yggdbhWIGW+REVC94wS4zI2R715l7eE2khcr8qmrGVSzgyryplVsENW3y14Y/u
Gzx7M60anPhc58ChitP8n7bpZeS29fI4jjfljgFm462luaKjLDSwXjseeImV1jM5TH1lyZIMg8ZG
hdFSf1js6b6Hcr7vapjVTEhL0DwCn7EKbLZXUH7Dj5aubcNwT+DDg4J0d3pcNM+hoSRj31xxS26t
XPgQAQP93IQunCsHQANQCVkq/ln2ST13Ednxvrv5dmGICp+mbt5oEtlfik6tt0e2BIwIlzpmlhf0
VA3cFgQ6q3OJe1uFQbEAHiYlMtBRnh5tDNNDBVYHabUEslXN+sWrirjEKJR4TMkh6EaG7T5xfafX
3brsdSnUH1S+M1AocJ6hK8VUeTMiYoJg3UY9b5C40Rcinf1tT0hIvruAVKiYoF9N3MbSjJicRry1
AsAYYRTxuTcGPIOzehwNPlWSZ6Kf7jUddOZ2vLf/jcjPXz/hYEt0o50B81n0zJ/eT5PCdyo01MmN
+7foOSJip1WHXtNwmZM67Nx36wiJBR3u5r9L8nxFW35d6TBavqX6ZL3NPtbkqjk6TwaXCg9zL0Ma
oWvAlqjKJ6qCAyFBv/75zSvdzSxxwHa+qEf6BRBLkS/42vJ6DdB6M1G1NKjR/lbJq7qfPaGiYc+Z
sqiAFb8mb/9l8bYzS5rVD9rEaFnCqCYCcVWZGRfHGkFbn+U5qPgqrvNfjVo2k6Tonbx3OOcyBgfX
X7MuLJrcfh4lCUlkPOYY191prUZg9ayVYtUUWh91U/dUyI+mdzdfOg/YTl9t8gp5L5xJGcAYCmsy
E7yxnbY2bbjyElexl5PyUnrovCPp97PUZc2iLUTq6MBSllK1qc67+BPIq/xGrJsqH8WS3MuAilZY
6XPvz6PdJosjw/dmuM9DrNE9tM/KhJ3vMvz8ar7h17t6jT33debyJ4JJ/2ivyQh/zBBwcnCPiOZ8
c2xim+abKs1f9gthpG+LLO+9soVoLAsghuTwMIzCgYop71giA/KCpSO2s8kkgtm6hJVLoitXNAiz
wXyxGo0fDfeqETRZPd5Mt4TJuJ/7TDd6BAHCnumr6dpZcupjOVaz/FRxHsRhiuDkG+feckzjR3Kk
qpggDDOott/pZO1MszyuuypHolGQS5wtqUymQ27L6H7ywDeM54nLTuLhwi0HAK4uTX8xTQhiStVL
cXsq2mFH2KORSORXT/9Gr/tKREDHYxrZVhAAC/Xy8qDQesbsYxFxC7ZdXyl2OmG2PVpYTTVIlYMH
s5If6OD8SWsyOYBpJDyqgjiRj4vVH++TTNZZh5Gr9ffqoTiIjhbAaQFOap6dTKqcEAf3YelAsSSr
FMvoFLAfPaFhaKvuf/friG/KkInd/JH4sY3jEkCOEvz8cEATySoKELe2R5pbxCLKHUp97bHARkGA
MFHDapc97nQm7u85IjZaf116vaHFpIh0bWnn2XwGOJ6oVP/rhFJUh+luY92Gjfs4T62biMJ/v13b
Wo2BRl5TUXNbjRXzjl8YLwkX4M47B8Xdb7JIXyBNpmGDDi8Ijn9ogbRlb0CDPBnSRk9rAIyoCjCZ
0V5vA/wLDeYYi//EUov4cUB6HEMbzgTE67/ld+25N0Ikay3tE0sFius6pNZMIfdgKNrG0GPPMKCR
WO9decqfkMoZC40cxVzQ7GXb+uTaAO0wYIsmQ2sB19U+58TaMYZBzShA2Jqfoc5u8NeJjhVhC9Ee
Z5FJ+WZ7uI53IM+B3gkBRp6sx6FwEF2YQRGRf1UxbJrJhPTI104D3iE/fCy/H9tlImtMyKLpW/Ni
uDxV5MGVHu5A55Ys3XVnM3iP1m62WVS7SBCFWQC9MvVklGbyyhb8P5aSfTpQlK/rZ37oX3ffaSIe
pgDg/fXjB88GChQm2M435Yt5gHvim1QpgOTNm5AUeCuZDifuZY+n8t9bUfvuAN3lk6rNhluVDSlK
NYtkiaCKokRGLjsf9IXb+qVQ9zgRJL9dWWOmFoVyjn07s6y1PLJSD2liW34I9k8qMUcfOE4BPoka
DrigcdmFtfLP8nzTCVnrL+pZR1DPikmCu3QMb9JWFYI6DnnakkPAr/sZWoVTQrvA7eoaztUHXqZD
t+LmuheH2jLibigKM+oahBhPMzorVkQw8Qzfc3SS098TO0oRJCR0AxtwLy+zcco5kU9Mn9qCT4qK
YUfd868/iDluMQHMFeLQ8Fu79FsuNWiNC7l3HVmLjf/3mWINnHoFhqDXTPr9PQ77zVFupmrUILuI
ulFKyHufmBuqiEhaX8N58N99CIpLFtzeof18VU2ns8vbUcVFXPSPKJy8SIfdL91u3bel1EU3Baf0
1nFXi30/Vsfv0lIH0+0KnBUyy+EqB+dkOnMxacmAOVKqJq5PEcIq+52qI/OlfcpTsG6m9RiQjmFe
tboCFLjcmjHkgbXbngv4EmEUZqbX60pUXReGYJk9RB4EM0XZ16bD0WWi9cvASLFJGTYpdlNpf/Ss
nndybrMCfsHc70rQFnbkOCRQB2g3BTIzg5+mRfTWVYbnm4Xne0ghh6a3E1dDO8ffGjcELibKV5bX
rHC32CHu5qQQONydVFzWJx+oYhrjbTaL8FjVW9kIDQh/jY7KN/J3qO6QmAduYId+gXhJPOPVKsVa
sJaVYkKSO21PoD2EKntmfoHS9D4nhTRt3DTVU9xre6QVF3v6GeXIkf5AKUVToz5Gkr5PYzysNka1
qkIAsZh4cdDPsY49kg3BlzZt8quMwqYCJ19Bd176WA++l0vO3q0r/2VvhPyu7Yi2vUrPKHV63U6+
+chBOwcDa6KiPVw7Jec39gLWtjlUN6YZBt1PsYt9+jasqRA7hSnqKU2ZbCYHVOLRAfuh2MZTL2Rk
xSWMb77pf/e8O2o5Xei6dxKsGf5lPLMvGr3gYpl0p5Jivsm9q2EwmY/qtG4setFrbIjitBDp7XjE
PRwmNQkLtshdu6/Cr0eJR3s3/VSL21m1Ib4+q4hF7jHuqkXl2/zyX8IYZS42pCHLRCG6Wx92UZi5
jMIJsjsV34rQjXAe8v88vSkIkUY2Nut2ZnBkudOsnSSWOT2RrOdTtEjHurcEr0AP8S4RqUtwYkYs
bOvlW3uJJ913DNkhwO0R4ecivONrPlZpeJaCuTmt3jJSqgWxzg/Gw8BLyc2kOYspANYVbaCRrpKv
wlryD1QAVGP4900XIUri2ZAvKU9VJSrl/4uuXm4yEvrAFZuQqRqSpO6Ium3v18eIp0E6/RmndJFh
a/rZQFCbZ2n6G+aJFwtI94XpXVVbNvYzbqhjnRhHwa00/nyiBtglRxY9JWxmIcsXRKAmyoCzDAWr
qItf+eARkXSSOQzrvghY9kl+47Om26eqfa94ZCV17fS/9t9L0xGWu2MoHoThu9ZuuvEw3Md1CNLO
kGrA9pYtV3gUruGjVO2vjkxk0hD1NIxJChl5xFVNmrpCjWV5u+ZXguqCA2ot3JB9LWZHw5sYd4Lc
K5EfOMphwCtjJwCG81CcJHOWqi/0Wu/Mm40WtgLxi23k8R0I8B6eM+0/a379cymaEe6KSJNl7LPn
ynqZ5+S0vSvTktoTZrVkJUbYpo5es+4rjeKpxos0wmXGcY9X57hvdCEGlNb97N2igf0GTqBbClwA
ypbeh2Z+/bV7HoUpBGuB7yMZl8/H5jVqXD3eRxr4hPFIQJHqpSShh4yqdEb8IkQRdTIoz5KMCDAe
xyKvGKroZ8VS9+5xZvDFJT9HX/DUa90UdOnzw5htwrgSuvulXq+gAqWIXQg9Fn+BqCfF62ZzsD5h
c+Ir8t0Uhe53v1H23PkgnbCc6MWTi//5xUiESLN97f8KLM36FTp+aNz9qvOuVUoPhC5BVO/fULZv
PEFhhGeT9UWoEhq9Fx/qLv5aULDrv2jKx2FZTVjmDZv2Yoo+5eaInHL2uTRNX2TeNTJHLsl6MwyG
BTq1rTmEPl2R7exL9iaOlUQ11TYLh5zgTb6vL6bltC244KfclhgwshwzCZhfgMBx3ceIS+cxnype
O5WmA+cNktbUbn5F8eyIcD/JjowJjjSx1XLwwjj5pZ2GAIqREgIH8XyGH9A1IEtJsev82KKgV+Dd
+5Of0BO1Wrr5dhDdylX72EIZMhkEOfScyflk6WjthqEuPMwT7dQ9HKDrJKLIfmclpfnL025521wG
KjPPOvg58+WbqjFvKSleApve6r2Biooe81m+ap2e/8X4uwTIKQmt6a3dDts1nOHFUTveRzeGROuf
16p/7zETFueRUhm3xhlqoJLTjNQBcCWXqt7DlmZ26seJX/2QymQKwkQGkSskk2zxtCh7zQ9yHqiW
FqR5JAED3hw+e5Ox5mM6CMz5ECmJ1e4d6DrwS0mzIjKEcvFI8acmJh+MgOozB85a+yrc1ETjaugR
veYO8vvbAiV3Aig3Ev73rhIQ65BIf2PfrgPHCMFEfXFX5bxgefsN2rZM2YDILHrSmrhheWNPe+AW
RVZJqboVmF7/Wb2hTI7H8D5j1Teq7sysSAph8WFM+xKCNpQkpON690yVDTzFpD3mfrxCoD8hFki9
KvmlbrcJqLuFUzJskzImauW+jbbcwS8GYcZSFG9a1IcWs2IYwzOaN/ysQZBNe8B6Cw2QUEsIZ5jX
FlGGuGFPx6C62Axvzf5vp9dKyvQy+qTjZdOw85Sio7S5idM0vhX6Ui1f0WnrNU1cYhOw9Mv7QmF5
BHIQp6574gnBpmV0o1FtIR7UgSB2gq+oBuTaprKlthwz+I0USxmtv8/6MgqSfVECTCeHzDI9R19T
8azmH1t7DbyaeKD5Dxfq7tMIJlt468oHyfA/28zgPfsR74yY8yq6H3IYdQH3VC0llRDMceVHGMkd
j5O9Wkzh+rgwkDwQMgWyP7ZfGNdweASbYZEgSbclD+SqUc3Ej5O1F6wlniq8o5xje8jm2mUDeyzA
c6quFGjCBlr/ByBMfYWRe9firzEbSgJOU7LXx/QZ6XDf+bljjNZw7sh6SWspo6nIo15UREvMXBLA
VW5FbqfIsPL5i057DwTwwBBkeXRKBeQFIeEG7oZt056gQm0Pn8TjP9vVqjzUlkRv89BiuWxeT1hP
woKodzj3/GabqgP+LJ1faQW0aKUXzRbNq2ru9eLzkdRpH4aDoJ/j5h8xo6h/evbN6bpaP8qav9M4
69OhZYUVEe2YpBECo50VMuqYRIemyjMHCvEj5T7RKP2t+8dpqINYoGAosTYmXHmZyqixSri3KBbK
f1sPA/rVb5aqUsTydBwkuLCF+DzSsolUim4j+HYeo7BiPsJjy7gBpWCujHiEnF2oZ91jDdWW/a0C
1coQPKNaXK/ORGzGemv//i/GCm0n0g5JgfsRVzKRfk6+HABLZYy0IaXSviFQ+x6W99WykQErDEqY
t/foJPhviz4jZL2RqAs58JdlLPFQnn+as3jCJ7C19YjLNcSlPV1vdWfOqR0X2E41bNCmXIRnCkzT
87PI9Dx9pM4N4erTu9YFWA96UjxGW6w23QUZYjf/3/leUVtJMmcVnHMiZzH5/nY7bRG4XsYoeIQe
GWMMi/eJ2kXYq91cHKUwENTZYiMyA19N4zJFm0qv/UkTjtXhsnP2ONF0EOk1E/UKqZctm7aTcMot
kJNjH9CeNiAUsOLZL5if98+4losI+nT+aLBeO5/CwMzEFYWSxy2rMt+yUjEphwpN8rjFlO1tNPn5
1yuL6Caj8PNt0F7P3mD4Vsxtcc1acfAWGCiEHfIwtFAQ5FT+pbTMU4ASiX+EU1v8wso+vePuCwLD
IwxUHiB4VkPLw8eP1vgiCIo5T8yFDpmaSYNyl4mLm+tlpa9nFWUJR2zLb62q6FC2qjgNBs8a8UtW
HKeZ60NDJ8jhe0zoIJYbgjEunTHq3crOTvDg3VDH3ae9u1Mop9x9/axlpN5nhlH7Bud3AJu6TzEj
N2GdWFHWPXCYVNjE/jrG9HFxHOj5ty9WksvO4oGepPmYAInzXint8w81FObLpd+GCquvXiwnW1b2
KQB4wdLDbBzDe8IJPcyat+pRWYg6V7npnNiM8y0rP7RIP8GiOez2EDnkuWr0G86DIyKuGwubV6RR
cZGO4HI2mC0Sngc8+ZqdbyJ6kklnDpt2tpI/pNQq+5A2CGnAAfz84eveddEdFd4jsuJrvmYEx0Md
9znB+9oTFfAvtNibAD/ep6tiDu3wzxPWFaSwbpesrD6aVojKmdy0iZ+sJBUOeClKm9qoV/yXBHuB
qcO8Jzi1/668Eb2XFw7MzW4ZZq+loVVJKzfbOBMJ6oMILAFtfjuCi5WswnudBnRpfe2QLTTylSu0
eRqwEVpGYj+NHaI69Zh6dTiVnieFS0zo0kjI2Rd1aw8d2TH8+BwXmW6qAMxI6lwhr4Q7HxUFDeQc
Y9GLwS53r9gch7TXhYO8OiMPpDIB2qETl4JOIySs2TL/3LGrrYSza7nTvUT/z7M/ph81ZvkVFv6i
LcoHlFKe9xeWkcJrreni5HC+qu8RWHmdWGf75owqy42rCst5LEXyA3wZloA+LNzYsj3vEmaB+pya
9VSPAkZt+/hIOZK4mjZDEQPK0FAaTPhSHwCulWVCoStSxMRnUSwSgH0WXflfl7ireEmkRXEeuhlT
4vIbBna6VC1KLBl3Pgg5gEhM1st2i/tsDYrYBBoc4u4/NEwdADmCuIV3gC0+yGyc0DWBtPgb7VVt
/uUntTk3eWttAqNvoWBTYyPkD78El0YdLa6wwBJUGLuB4LLtTgGdJUASK271iJdYHLdB2yQ7ynPG
e1/pELF3OVhdrJKFT23EWwSKcxdqqn28xJdNJr/+dvlxCkr13tyZMGXX0sgyYaQQcnDPvR0oUCOe
BEgq8ycoQwZ9jT0dfZlEAZBNv8+pabfl+cb7FPPto9UvSo3R/Q3UUMWWEV8az6dgniDE2G43+gnG
7T7SCuDd2bA8+OZERK3YnS1Xz2cnoj3cGet9Ut0KteCE3GF9rQ9h+EGAAYZIxBRajfK6L+W9939i
NSM6stwayqI8JTeKgWQUTVQbSsmRiR4Y9xvGasj0oYYGOXSCNHyjNgOwqkiOpdRpLTQKR6IiJqRf
nWKMSVf9NExwqHnORLePp6lkPDxOzBvRlXq66sIggy1gfYlnIqTpbTclE+0Gh3fN/3GGU6qHYOfR
xKWwnMPYF4w7+oYCOwq/sYhxNHy+E9g0/xUiIgBuBtsirKNvrjS2j0ll5Eg9+6G4zkMXbHwofOlL
5Hbufc4Ge7rlM4P0QlZmWJh8uzyOcD/iFzL30yaUQzkh4yB+imnw/3tyhB9kRxUuUFwbQZ5dtT8b
piQT9E4KPXW3icKEYgxvPyIDsCPdJYZLnKeRa8glDNQICpkiK/ETOV1PS0IW0g0d1SscTcN5oZxQ
0YBrwtWvaIux+DuZ9XkT0tKD3rNXjPyE+WsKBcpw58DoRcqBt6YvGRKsf5b+BLG9QHuGpND6wUUA
6CsWIdWTFIoasEAWgDkqSJdvx52f4b2JbOcQCrxn8/7wJ8qUi5NvToChb3V97kelEt34OGh8JyKF
RgSLvoYjfo9MqFMhxB7MtRrFlMEi7ROMYJtJVQ9K53OsC1dpFe027Q0uLmLvcm3EY9i/gn8wydW8
F2J9niLr7Y0khVMvHrDOoPEUX3llV8OXjJL7VTfLKXtDDLS/87lt19xDF3JKpdpgfbp6GRoJmdL4
19DocsUszaYwMtdZTpoeKbuISh2XDpNBa98GdYBW/sNaSqktq/qPkmBylAFgCGsDTDsO4dLL+OqF
VQhzquBincu9+4gMy7+C3TtrLDedWScHkYpKZKfLzDByxJtMTQ933IbGUv9Z7iR8+ToyunRJko/n
RiQR8Ni4j7+K3Sg/EX/LhS2m92RiC8dzU3ZmtkpOBSzImDvM5gL7YXtPePvlRI8i2DVcimM2yJwA
O8U533Zq4GaAGSGYyOCiVW0Vuf24Sy7lsscu1ZTbml477jfBvVazXAnl2uBiMho1mxxhiH8cMLOL
QUIJmjJoPm7MV6HgQRimAwX3Yml+cM6/9d3xGz5ddEMuG8quIsIm7fZawEhJaEK1/rtkvcWksTD8
zjj+oVU+QG3an2znCh3/FxPri3d/3GnEJfE6KMgpji+AcWaEeXrX3qJQ5kiMGgIIy5IygbAAO+uj
ti5w6spACStcEtkmwJR4uPeXLS70MMKgVuvozH9TCG4XJBtlDgEgd06Cj2sL8VShfozKTOwxFI6V
irVCh+kCotm30dzgnEpzArYGuWPRXjXQMjTMWQUyfgmwuk6tzhh8HWz/dRyQXfNmqMGU8NdYTD19
UsKHxh1+zfElw3MhcoCpyt8Ey2Atb1t01dm6T9Nk5OWc4fgMgYhNeu+6N7g4jKQrhGbcUxJVJ5vG
JaWu1gbsGdkukSZ+WfbCyiL25Nzl3brafoiJd2kBF6f/yYC8bFW0577ZCtnzsCPIOW7UAy6yT8/h
DG1NWM3OjD2BTYkw3VWn36bwY5RYKNFiLnPTvRPZeMMv9NLSGi0MSYWE2fBSzRpNqD8t6JmWe1qN
O5c3PIGFE+0ivjrcFbVVI8eBRbftVouNv69TXo/Xd6Nq+uqBg4sVquqFFQ95hCmPzHZcB6uBEi1F
yDuShQKgrGS+7UlwOa0alJUI76IFP8kD85zWkOXI3XPxsPgf7Ywz3tCcfGXSRXXu5Au2FeK8wf/B
bMSQn+3tfMgH2dUz9U0Cj8uoX1R+tl9veQ++rrRbJZz3u0L63TulT6NLnZtkCobquVy6S0LrrGAQ
RNbdqxajnrFQcK/PDjvivipZBpNpiJMFUb9uyIbpSPrbF8mpiNSEC695K5dJHhr3KQtAwc/Uwf41
QxKZARMLWjgWnbYQ8/CtC37F9SegVYwSLtTqXhdKp+2lsymbCOG5z1ZvtceT2nim36AELifV3ZRv
cNHmF7lat6JlwLwbP86dT/lYk3MDLMfUd2E7i/miS6IyDyv3n0HkmNZ6RF6i/NDOZ3Ljy5gAT9GH
wnCTcHwcY7AYPQeCSXvLZ51wfk9i6A9vOTVHfG5pHdQl1zKL+QKAW6WKyF+j1ixVC1pmqYj3IJ9U
hvRBqiNt5OUnJCbYGVqwRzjnHHQbHGluv/dj6exvbayjMdnC3/WKGrunvcRg7CYSPMls6gHsCTBx
tsTnWLLWsjuWdkskYYZQvvbALKXbV9taYPpK5xOTdBP5YOSoWTw9/l18oWAXVPc7ayV4xMKMdJdn
4UIa0nhGLPUma2U2eeNey6Zwocww7sdaP/dBVlTcfgVcFDx2KreAx1afC4ejYkah500H5J64RCzP
43amotPkQq9Smj3w6SYnWcwaErIu4209Z7cBuDD7gWStuNxo3HWjHXjkMgBva97iQ3b789fybey+
L53vT1dwSo/gA/V+eOffxJby8grMW+/GItyrDFJ4P2+vpe1PcHgCBWbjZnjpvTyeB4msw8GMaIEc
6OKQ22q9WlMjD0PyMVe8rXHdJ94jjFnsmoctHbqgqJwjPFLqnVZ3/4Dgddzhi5GkzUltUO7+egaM
gMhfFDlpwS5zB6eiAimtLe/ICwmcGSiXmj7rgQrIbVPRUl/utT+SSPdDzriL6NSAsNH11LFuGxTb
vM11EGYCYRf4/x74bnThJ5rGthwy3QO8as0xiq1MjJuWtEw5q2wF352xnPL5YrPewk5l+hKyRA0E
zeRPvDmK0wdocd7I9MZ1JZaN5gx47pF2pnu/doLXYZoMMbvemDBbBlkAJF5gnlil1QG47ajUJndK
wDSiPY3oC/4CWYnZt7w17JUJ0LJ0/5HDN2+lQeCv3WLZ4o+j+VNv0h0+jmRiFmhJFLEtWJlyR/78
Amhg+7sRWowkvZHoyynuvDP2pYuQgXrrlb+wCx0O8V608zqDeNztuDhz3wLLUUzHkaPDvLGH6+2C
afilSsy/Ri7FV+S1B+o+aUkDdiiPR6nA5crFZ8isOxPN0MwBGZuRb4KPSiMEgfP5ioD99bz7Wn5y
Gu5IHI942A5kEvYul/7FSdnevRpsyQoi52/h3ZKQq2ZmG6qQ10GZE7xUSqU7fCHR7RYL7DLyc+Ve
M4FLq1rJKvz3nUuCXnGFAAi/9yQePVExYK8Brx3sPqYZYiJLID4KXsSoubHVW5wpw/qsfBeJRsSe
zcAt7eJ4x9FOBKf1nclDfHIgKAzai2fpJOZ4N02jZ0EofjuVtjCaCZmH2PaGwEkibnnoOcdPSpN2
3LGJT3VlhfaT9Z3jMRjr/G2KxZcdm6hGI3iCYgZX/qPxw2P+rLFb0NjK7jXZmT04HI6NYdbwv/q0
Ioi2e0MAVKkx5xEYaY4MMNn85gC66nHWvzbeDQm/IV1yTtL3u60KGofLjWbCYzqvQyhh6RSnmom4
EmJT8oMd/LGsWZupQTPFzycvZib9moEO4x3xKcu5jOTSxYFGcx7IjqBeF+fVJvbTMYVCpB+4exf3
zENpAfGuQGxMiT6s/QV/SCThmFoD59lfg1KOtzo3EwRG0HVhR5uJk5w+HsPIZXI3iPEsNhbvRX2M
nYzQDs5pJ7yy+gIT4WdLTOQhkbPeG9p10FvjJCbuG3r0SvMHMqT/AjzOiCvPSMxKDJKmELjyvN0g
0DDN2GAcmSjWNRBY0B4FZXaKAPFmR6c0Lvk2hLFFpZ4JEvi+k/QRTWa+XgInuHcMarg8/ZeiNf+E
6eAHOBU7aYwZX4P6M85ewA3wPrBZss8nBynLR1G830FEgnLJAvLOzcsT7my3f2Q1x0wyzbEfucV0
MRd4aYaYA2h0Wn7DEKWzIdawPE+Yve0xpMSk0wXB7guty24ryH53kXgVkQnWmJsV9ivUMWB+rkTQ
XhL+P5YCeci+bnP2+C3Aj4aoi7YFSQ+6R+b51fFQmiSbEdIZ+nQ+Qg3CJywgSsWXi3gPodedgerp
+8hsAKLbcFTb0HfSuTTUjvQeSMIKesl+qXk9NXvj5ya3DWfMeLvnCjXpkBFa8Tz53MqfJ+cpnVbS
dfkgPT8mCfWNcP738DerbddxiNV4eGogZs92JZsJsgrFVutjvI62qBn8tV/eO2E/ZAF2MaLRXbuQ
Bhmijzvo4B1z3VT7tO8hysuqnnoqWheul0Dg5dT2WgX9ed300jtYjyBCrf/TOxZSc5NCBPu9Jt0a
cHPS/yc94VnSRIXQ/81rHWz73rrVtGCrqAwo2p+CJnuNbfFRRrNoOXb2eooooM4dXkW29TTXz0zC
ertsFYGTVvWqL1+oK173TLbiRViCnVa6hsX7+3rgfsCzSlY5wUiVBBKYanl5OLxgwMH+qNRdGIh1
wlZpT4QeD5TxMtuY0Wr5ox5QqGaBS0shkMpxIrsP8+1Kf45tRteKznhNj2XEqNB1diJ6CFSv+bHg
6Q9pJYgoZckRyXlbF6Xtpmq9PWW3uQu9SkGNVs2Mj++XTlH4AqRQ4I8Ba5ljeUVy+Cko323WQEL+
hm6XxgPHRFOQl9IsxoJRJpOke3B5c6at087S8kb/Id6ajyKiDXclqJGspaUwyv3lWxFxGo9ps1gi
Cg1X/QZG0kwym2zHUxnPPgqS4PAUqBH/xJUlR3FENbVrDF/whF1K1nvdOleEuUaTjguDVHASZOxh
LcS9YjP2hC9FNO2bqkkrim1a/pDNWZfzItZF4k/JDJfut/gN6fuNqdbQTH3d3RMKyIjMoHtmorjH
S0IROG0JTaRXQUB7V3CPc33uN78RCd+kN4RWvDw/rHzfIbnwl+s/PT/oDCjRfOzLLucZ8IkYvpVK
o5IsPZkUAlo9dQhVGZWepSJClMi4AXGpuWj33ULqAR0erGlLA1ZXrffdXFNO9ocU+5lFBzd7BE6e
Cv8jpzQ/ORcc+QOt0t9bAvLn9J0hEuMwpeKRWBYuKI5OVTbojT9jD7p6sm37tg8hIZDTXk+CYTRR
uPah/40h3rZHVtDgHyYMTsAZc0Q+5OWDYi7yFwzVadtvUCkCnQdUO2o4tNGrftFZiHB9tMHBw+G8
6SmDlwZnXobY7MtQrowxHBJc9+epn8ij8tMHwWb7GDPFgABHgE/rSqSyD5La6KtxGZOgXiyqsA+k
sYyr9lvUz7ITcskYP5EzW1F+fhtm4cA7PtT0z+WYGAKjXquF+qv41zLvg65ZSlDKL84RGNpczpW1
hWBb/BALepzeWj79YPFlSJ3J+00kS8cgdKLUTe792j7WHKUYxPcT6koa0widGO5yw9Dyx+OaG1op
k1F5T9mHxZgZfxs0WJOeD3tG/2svu/smtj7u3Axykm5LdDWkEc3EsmxXFqwPwRm77acPfvfK3HMs
HzOmimckL/+gMEk/Hq5RBX423o2+ttKwsqzQSizQhXZFRjG/CepErkBJAlwOHxwJxAQkJ3sQ8dAI
4D714mR3aEx3tC7HVmUKTldbF0OwkUWToErX8J79jX23mCC/E0iWUk6YvuwQhTUaiI/Vwy4XSnz4
X0SbqbGjX5vJBVu2dZvsrR/5p9Aiveu9KrNZfQED0ZktLRiKgNAXERBd04UVvJekCgz4HQ9xZrnI
fj/uPKx80+gtHQ/iwFS3ByIzjKzD3xlA/yx+fznPmDqJyqzpyztVFDIySlYFKj0iofNLrCWTqNPZ
eCxqKXkjYhhpSQAwM8waKPqVKEXEY41eqVtzfEB1s6Vpyopsq9BEEBXQ3OZmzWhWJewIW0WxvqXa
vhb75BdIlmrfcIANAFlGCV/i3RtruoDEhLtQoOmqDMkK3Z55pYF7CBeaes90O8tSnIh2euBV1hyj
2NJlO2X4KEKdYxGz4Amh0H3j0cZ0nSiUi2IaZkxR7CRSl+LE0Q+URe1nvuLtHnbzC8IC+vbO97WN
PZYLRYshvRvlJ4wK5WbdYaag2NXyWmLsgwxbSAlkRsFJ07Qq9wvBE9gDALIsG8wRcfNvfK3ojjjv
FSV+hvqNqFHq1XKgRKG4iC8IGHYVJ9FRCAMkXS6tVlvZk4c2YwzanyaIEuEAo+1s86UQ7+tWAidp
0exFdv8P8NxXVT0V9oGaerf/8STL0LI12+hFYW23yiMULawK9CT5Um5lS0PVoHe8BxUKjlaxhFmq
3/JMN8QDfCT8T3qkXyRsfn9Ns+08x5xlVi+ixv28+mkdB3qFnX9s5BDI9FrAZVH6NDaXLSwRla9R
DPXAQXjhEKRkpX13JOdU6VfnSOFiFmNDoC2jJVi4aLZO+T99YvukfYMC/yd0LqSJyj04GkGdnwgk
02OBFXlRcq2fvWznkKfxWaTnOhLMkibcuL0j14OX9z1drM0grU5BMxbXxT82pTYat6d8K7Fc6Rju
Tj4pi6d1cdIgSyA7SGqgPtCYbFp/iB3Y/2SU2tThvq9TTOCdnSmo4sKd3TBmfjzqOokr9penBYhC
L90UoJrs9LTKzd8NJMnUCBBJYRvePwFKaDraSjCqtFp8wiV9Zdxfw0/ZbeNaBwlA3ejw/F8qD3Un
sy0L9Oo1NegjDqAefIWwMfiFIWOFHeaMPvOOii15JPVmXNIhqdqWRXi0IY1NWXM1sFZQ0xp40dsb
DPLewKFg9G3Up22c+hOlTyrDRxXyR43KamRwjlEI728mRo6GdPY7eo30Hh5m8yxeAyLo38AGzypu
9yqzWmsONOvX/6jCd2GtWFty0UnkBf/hhwMYUTkmDfHIeVINOmpXOQyVK3cHDc5JMsPujnhKHdKJ
qh2KHJkiObBHeA0pWzwefAz+YMjzvM0PCO5u9Dm8eYDZAkcA2DhdJa6bx9HwEV4PbGfArT4xIUf7
8paRKl+kIHx9mvaqfaPo0BWHbuoHrmrrXYYunUCrXZ6cYMmDuBARbYj4fTEw21jvD3AR4kXuEyiw
y3jYgRh+1JnnJIThlbPzl3cxQlvLq0UffcR2vBv2o2Tbik2s98dSgqc4F9qRv8zSzBWiEwsotIQS
/2PZ9frsSUQmnMyYx0VzKZpw0iGXGnLNgpf1oIJIFTNu8r885CLRoYaI6T2FX+6X8dv2o+piVzi3
zXQp4txaj0RcRjT1pjkZDWwsAyddB22DS5CdMokS0ULB894ATENlfoHCd27hzyjWVXqqDYN5ffle
nhQwlqqbA8tFQTgYBPXMVsZuTea3dVAULKrjVR6uktBj2kUbRJ0Yrprjjptr6NH2+aEAqf+jVejo
JbSwEV9bvDpNF0z2PANY8p4Clt15rpJIjIDpxVvxKtNBFS26O5LQpelA0OctuqzDtTf1trWnY5pN
328iYa4ymZmQQsIDBOmyoQCLdSPibtMxLwBRjkUycWXaJH9uQtFrb8xmTyVGDiAd6dFRIITvHYvc
bI5ACRYW9Ao1X37TZcOA/iL1dj5/OYBffTMAwG4b/kB4hjvwDttSiQROcYKT5z1+GZKmNdahPj5U
EXXeVIyT3YhRIJBKNLCClxIM7VhJh/uSHa8w+t7UbVRZgGyw/dchd6bbHZjkK0LpmzWdnNnRUL1h
XW503XZLm+qhtoQwiooRm/tHrD0O+XeJ9KbOjNSesCLmWs+HFhmG8EdsUEWKnPCtR3rxzJVAC23O
Z0zStiN9S++eY4m2iLjHEoOQM+ZAwzHi+b0XJS+2/X5VpWwRPl/0jRe84Ky96h6qI6sB8YZR+VI+
lfUeIhekCO8KP0KlIF14w2RAgubK9WGgt/jp7xtk14NmI62toJMvZTcT3SuifSty4HYfi2iO+Kei
37h8/NhywIrgXfEbxnLk9FvTM9XgqML4SdZRA3cyLAsbXKlVkFne4gApC7GMy/F41l/jJs8RKVOr
6yZCaqFLl34V+g4fQJgpRbz/KmcvwzPv5P83422KpDH3asQ9mVX1ZgjkYpoRiHqxIWxL/jmHwNug
NCUIrKyAzyOsM+5leSzU/vsxAhGbISV2LIk5NALkvTibB5Q1vyIGh3To1jqgqz+sbIzGP4OKaswb
ZKeUf1p6EKysW5e3nmaACtsK+ouABd+M3oZ3ukuZkEy6/wQD28HnvpIJ1wP8jF+aLFfx/dY/r9bD
Zp7jlRVg+j7QkQKMkaPwOP6Mh5G8QdFD3AE/KL9O/WT6GNXhv7BzIQLF4wpRRnZ5FwQggkyD5Mty
UIgMjktZpq/V/tx6lAo368fyD/4puVXbhatPJ7l2AyFouiYAClJ2XtjY+54WEVtYh+pcjYWXMfqz
p9EbXu0Ong26p5sQ8rY1EHpPu4B1pED7x56v4AndugT4CDPhTN5kjMfxJjhcFzul/ZLgrUfbu8Gq
Uhw3f9VzP23CraQ+4PTGguYiE6gfGb3krn4oTlDbvGGzj+xF0b8971UBHehEx84NQYppLprOVRpe
4N2zyA6o5tlVGG3ADsxYtcF85typa+icETwgM/WOg1K8DGdrTULoy4iLOVs87D+xNbuVDiOSN+rD
TRCWkYWPpgNllypPWXeUC+JeX0mK2XS9i3KnhMvwraiWWYsSHNJpUA8WM/xozqH8vi1At9FpuNH3
vvXpplFHF+cFv8awEUMsvTQk+VuBrEeIiQvW62aOS1JxwQ2D2+MgfMnIfDuONNnP/HsKI94EeHE5
DZz1TA2zpTuN5En4YPyS3G+mIHiU11+FZg40+SvAQP/Gag81G01AJvOt5jW+AtrZ0eKuXhqeBY4Y
PLN8qXZQsn0LsfY6rzdV7Cf1heuostog4dkoO6VowJPkKQaXz6x1KKLBi3HVDzKSKOALV/fTEj68
kSi37NBo/UdJvbo1EFoIPYsA5UUdDTvpmcJymAhltym9fOWSApaYOxoed3iSomfp5//DY4/hESGb
G11VRUamx1BSgeZqXoLiuiETGWEqara8Y8Y6MNRy6qbPGwh7yH8L+wXgLhvL/Ni+hbU7H1+oNjtO
WpaS0D48yI6yU0cLmu+sxqBuYryE6v/GFvNJrEgtsUKO6nW3JcP2WqI1IATyQ+hDzoonV1v+B3fT
z5QaK/6p/nQtUFDQc2CwseODr+BkyCkZsP0v1q80gJnpIGS9l0iz2TTGMj0TjiGi2hYi5BdcR7Up
M7v9Q3LWQQQXQp8DKamyNJToC3Q/69DexBvJ4HrYCtYHungvO7NKTU6luNF+Ce2Is3OqJ9IeHlkz
3jytZOhV6MsDdrxs4xNogZDaQvlY/fIVmZTruBjGWNzYdJRwrWrRUZEx1dtTMdEICl/bm6aEU/Rw
YKbHr/WyhZB7RGGLpNwnle1TfZEg8uFJEBth7vTzSFaKWYdL4VPKYWBKAZHOSv8np/zHr5IXWEX4
z4KiVJMqn5UZckdllvO88D2oKtwP9S5O8NTIpydBI9oKcuTxgIua/1e0gjU+MQ6Dd1JHXN1+1lRU
e/huJQPgbeqW3uueShoCg3Ko0CzmYvMwu/GoUFkAkTlR41pngjcjY8c9PAyyJSOyxnpR/kkFrGiW
Y+GFiz5sYAFUkmT3OuoIuR+AjWHfFH3iC87NRvHVLcHaUdLrb6d4Y9JC7o8Jy21QiRpciVS67sGx
r5pOWbmgYX6kaZDJa92WnefdsynvE+lFrUut5er8XBbWkOiEZQPY+bFXR/4un2m15LLHdozAX4wy
5augFtJ+8jkclYIHVSUpqS6gDF76nv+UDyEHGkH4B2rlCe3SPSgRl3USiawi0lj2rW4/0wkKsPlr
c138jumc8gCfOKDOt2/Ue4a8QT4AGbnDY0dwCgSclgTdXOB1W7ZnlI2U1JhAa71m5eJ+O1pATIaO
eBRlqziaU5efaMN1m5VG2VcM4VryJDpIJdM9WoxMZrJ1AtZutR+jBG1FZacTKcTfFpYSN11XAqJS
glDAX5ubbo0lkhhrdB7B43mXNhrQuEGvxIHLIuSWojGaeE8QfjKNo0y1OkitLZxWv/t6LRJc8Z9b
51LOW8OEYTj1szWcpLzNPbt0RG7VeIjDqaGAhHMZxRTUwMoP1WzZYBKE1YZmiNRczwOiYDTzpxD+
utOsPSfDMMbHplFzND8B52zQPIxW0QeglZ322PrIKKhECaQ1yXpW0d+oAZY2pq1Lyslx3yGXVUQ9
1RBBThRpyph70KuQnKCAxa3HxYmuSzxUOFE2ssOZpIAbhc1wmRYy4x1JEQWq1IPZzlD7aarMmRJc
2t2+eCuoFcEc5jsZLBZBxxsi5+XqUDCBsx8Gdd+ejZdG92BK2Z/XgmSX2V/XjiDUTQZwMihcLwXE
HCOonNc+dncxaTlafGBB/AJvuAjOj2HY2FduLgUexPJHTkykHTlV+aJ8qJM1k29twrLd2ATlADnR
A13Jq/V4T4zr2SvC5S/Fwq0C8tzaU2eEVkeCMFjvKirafq6lTLf+EKq0X2+pAE9lSSTdJIX1D4Jt
UGyCjGwJJYiOtrmCPkKtzwpWiXjug1HWuRswuH0wxTEDhKIKVYfQh49KWqyIqMNXU5AknlOcWHxl
v4InxuoIZT7+zINKXji3aegQeOEzhV8jtjGMPa3eQy5z9TxMb/w0Zvk0GCyAADyqUU7MxWmrua+s
UTqkJW4lBSKCgFnM9KZg//QQoYSDLEsuLhETEjO/V5WFGMXCgfGx7Eah3JkcYFymGFNvLg4oKR8Z
RIIkeZhnpvf/fkxWqYADjulj11EBvidc302uNvPVfpUiWt+zpi34yAmT7C35A3Lp2xenOrFuNNBH
uGosiWAw0Dah7Xg5uHCLs5YsjD2APjR3d2wOQLZzllfDv4dQ33zTDXYJVW6xVpDrOoHk0EDe5W30
ly/Kbz57aycDJXODlZfGT6S08jZVJNvstdfvpnBZMv89v03hV9/hMBPr+epq+UJIW/e7oozEU6s1
ylE4UxXSzRcHtB16PScRapAnquW+0F+7wMAadvNEKFpCAM1CE/0pHi+Depf93tkwTGgHdVnDwGD1
MRX1UXeoXXZGcPmHkEC0+n1RSDIB0okS78avKdZK3vXcveSFZfntbrdnIfht1DgvRpTXpnAxGgTc
SBmC7yJEvReHpmgEyVhGVMJ/Y0YSl7tldwKiDZIVLNjCNbliK6swBNKDMdm0NFnnQIfTNWIwfwmL
b3xkLhqV82YK7DksLPqlozE35lHddsXDfDHoRhpDroOTnnP8IPvMbec+mec8bi80H2CE1wSNl9D3
FOCoDNIyOpAGeFelg1Yl3f6FIMK6bo5riKuIogOefc5cZFKugIP98fKT2EPdJE9sTtOo/5x1vAYZ
lvpAL58FuD9z2+C9diMFETdRIIu7kwMEYcofFTmmkC8bdrYURUg4nWD5C2pJdQuOHSe3JmKV7soP
eQPWj5Fv38D8n4Th4mvyYJVsnQSEqfVveB2uiCKdOAx0Vh4e7aJRp2W107sXxWklma57Sg4SxBAT
Bu+ZeBFwLWBI9KQlK5VkAh8ae4FcapJ+Wf9oFVMwU8WobciQug6NFsfX/AkFIIr6UfCZyQyZclTq
9DfwlMQa3LXGbDqiXvqP2YJtgiGKbHgeeVrBm9NZX6Kf5xPJQa+vo2V6O8Ysz7RDIKk92W7+WVKU
nXYA62O8r6JpdJUl+bPdZseVf9B9tZQ8NrT4QeXDwaYaaxxcMS+eHn6XeIi+7CM6eZgDrwA+Fb84
XTsMds58osqq9/XTOOgd5v+wlyuMK5C+eQ4nFuKPiQIcFtT274gnaYgkRq8yt6isQKsz38PhNla8
/0svegxj9oXExGSqMCXhBuayLKqXP2wdoOPC+Ozg2YPaD5GdteIiv0hubSL59FriSma6dLhwEuS1
amXHoqsU/UvxmPqBor0s7sAicHxOMder/g9QQ45uoVPcCx1/S4fT2v5rTBcKDS6l86oSi+OwEPJP
bJZIsIcABFTZ7LoL7rcHVaWxy9ZCg7jfx1bact39SMTcsUn5X9AOEQfSZ/5BhrnORNqHF0hc8heO
DHZZFmfM9CQXEsmVJWe9JNnZHuwj/OiepKcn/gUrng3jLl1me2x+vBF/T5Tma2TLYEwlHVG8V49W
9Ehz7N+6dTTPFuLFNgALDnCF0aYxjhXmLdqQmxGVmaXpPepVyVoW3CQYaH2Hb8AXysFtjmPZKLOa
NutcKYnFhLo284AVt2hPw3uK8ym9cSGdU92CFs+bMDtp9g5KaxF1Q82uahzp8+IjBLHrOTF0IyK4
9sHtX6y5zRdGkInMTwfvI9vSpNiAA4DrMBC2jnMmlKk7UKS2jksWEB96TyykkI3A2vqgMFlchNqD
2HZKmWoqyTgHtlJb6p9LpJnDyELqRlwiXREWWPjtrhAIDHwrwxv8LwcuI5vIC20wmDXrpHKhwWud
O73Sj2C7iNrOUDHxl6BftnzU0CxTQaPx8IWmpx33ZlOSHunLOKt21Ga6j8FJsgCj9GTnYTQGPBIL
u/+geTZbeBua36gaBZOStCkXhDPgNavy37t9AoGtj+s7AK5CQX4r3O6o9tG3fui7SbEfklIEzOm0
2ws3/ad0Ldn6ZoJaAdOiqbebMywvrbdhZXVmLZTETcVkVJqPlUnoaKFv6/00lfS8+hP8ks7JFQvH
FxK+zZm1oLOtyU4i2bpW+wAX3SIJlv48u/baMSpM7sJrPPGkTBPyRYit0C6yiUarvJCHj4WnOMi8
WNXSCcYrvYe3K0ehbWm+BCwGKtiGoZXoFv3mFtaGJxsFuhXHfXh5KD4SEgqt2odJwG36iTzarHOX
PkTTaDAoMTxUn67LeaiHiT77QSY5+JtOA242fiEpgmLNRqk+8PjUKGmFyG4J/Ea4cArLKAqzih5m
UGNt8dB0y2t4BhIBq7JoaNUcmffUnVaVN5+rAVZdlZVku0ZeMHFXRLKAcvOR2fghMmfc4moF0lTZ
O2l0APqMBBqFyjzRf0NL4ds0Ejm5dvpyeLnEMM9XqVKXRkRcuYcL8hZKcPiZk597nQaXsGS1VER4
d5+zKn8hQbLxQpfSckviH46dFB19b7ROLrWEkAKfNHc9eGuX9YyPGDeYRvXmCzP2PdKAWKnZ553R
Fw5anbMjG/YceLykJd4knSJ0nTtzwldgZrWHchjyPxHH3iYJIaIvldDLPDhnvFKXJnwevNhCus1F
ITtZqCojULv7RP505NILRINFzOfiAzX0nHeGaQ1Nh/QDiZMG5HC5G7NKExtGXB9bD+9Pl/5abepV
2JmdXCwtIhZQp/QVxjCpp19aQpfyms98J85gOuDj4toP2xk9BFB9V20UYQinIUN+CUtn2KObi6vq
s7B/bw6byfwjAS5Z39oQjcCrw/2KqnD+WTtn7PPYyGlrkT5JQI8wJ61TR2KB1zYy7yVjlw5uLnwn
3nsqhfiOCTPjKyJAiRHTRVajBR7TJqdx7VSXXx0+9whvWMAf0LET+I0gsVIDcIsnjDY55df11y54
LVmeEeWcGusaSqe2byJY41hf9co8Enenqc8YTGGTt2jRZS6vfI4Z9g1CUTJXL9JQZd+hulNmBrGv
9RJ7i+cOCucxsGxU0oXQu7oLI1y3jbbpl+a86lT8gAM9/1dUoKfdO2gPJe97GW0a27lrlKZ388xL
ULAqA14/iye8fopjnTgoS3fNfwaEaHxFPCqZj/EG1Yd1SG3/UrHEforUz3x0qTmEIv4jzLxnjkwC
vGVIg3MknsT/f7Cz9ZQl7AJYNJXlnN1mu5x9etkutDsbyjQbVNvv+rZwKoHvbLReqTR8Knd6sdpA
NQwhuuVFwKuUGs1e/tN5BLApFdHHk5m0dfUShLu04mrspLjZFj7kVlOeNIDErLR7G+knrtsn7Iyu
1MhD+WcNnveSstM2IOeoduo9LuQ3xGDlOPOCldrRiChRS0q6cJJHT3AloPdvAi+Dxx7ME2FZ32f1
zES2A20nXc+DCNVQuZ40uXsYmxZkZ8nlePR8SuR3OEfMCA4s0+batF9n1zC5TbOd5iQsshnLY6q9
Bs54PCrr7ioRrBflGbAUpPHDTOYWTkGLA2Y9Ry4pbAIbgihUnrPR+ZqSgCNLxYqkHGkoRBQQTQyL
1kihC2cOmTi3oRL/0PGDq/zaFmwHTR/8t8qhSU0hYf4UBXjVe6AaQ6YWHrbqebXIHm0rcC5OHnjz
VsUccIQ3ZeGREwUnesasBcVHE5m+xvW4g2JYlICgnQKSKikOMc9UZcj13yeCxieoARjcoQcO9L4o
rDtOcHaAEsZDQN7reGRws951N9sslODNlq6gTNsOx05WoPThJhbizXMkX0X+wy+jH4NzFv9KgT7b
gvuynDvuVAcWmg5lno3zkCW1XTXca8WLXqV0o1eItTodkdLwyYWtyo7rFrjVOjobWNhidHLBEjLo
I06NPldgznbLpKpAp9SkmJsK7AkA1ExZDrMLfW6/lRb++o3QkmylNBF0U2ZisnutrwrsGIccZOZy
yY1KguRQ2Hn5wCMTGpJ4IWLn4oIBEA0lKmKyDAfVjnr/rf/Ol9xZ7d7dwU0r95+r2rmvObjxCNm1
kVCjXGtHiFWwSuh25bKyva4/1PjUIBe5ThjJMswe44cZD/RGFy0M1ZSqjOVO8+X9NRWIuO9QK75i
5CSxEdy4VtX46aISdqtOFE2MbkOrgii56Y7cj4pA1Y3YHjqxiAWziMKeUI2l8UiD7nxIKhIXsN++
X1nPU0nuJJz/slP19a92iHyKUL11Z4UX6qOGGF3QNHNhcxKyUCNCcVSDWvKGOFfN5knNtA75KiBO
PYnC7ojble1EXtOYNzc73aZBwRErOb1VmHkwtrsHV+EcYkQunDA+nk7UkJW1RJHnWbnRWzWbL0Bw
wQQhMwepPTx80A8U8mlGpJamNhKIthEhKT9V6HB4MTTdTQpuzNlxI2I6b9gL6ptxw+HuzBlGCTOj
0hrx0uy86UeNq6DRSK2/G1nBPl/5q74pzttG8UnbbhfH2iZa23rdn63+5cKURfUjNpfc/0fScW5y
O5N3o38etKv7WIrvGnYhMGzVP2DzU+WbwLKJq/SYZtF4pjCoihJ2A0cBKn7Fal18b/IymbUPvrbK
HBNwKJ9oZ7aOA7sWaxNCZXVGYgoKuzJx4/JFlTNvRL0BUoyawV9RWqyg9Y3qJXg7ud2r4V7/ZM+r
s/dNP8+3C1F+4LverhDanI98mCwkhISW2hgc9hR/Qovu85Io6PzIOxkgmdzg70XWPDaPvUHmA6ZW
X63og1XqrtoFB9evLQnXFxJUglZnoeU7EUn1ObsSYRduF7p0I0YKH1IwAjSukUzARtqAswo/Isth
d27IMdiL0e/GWht1i/yDGP+yGryNqtTtzDYh+6eF8T32+poB0kPgV8Em5SLg6msAGgR3JCv2lkY4
DK4kYmND4suUatc4ZV+clgwfMmFIbcBEHF5JoJg53Uqsm+GlQwIyl9McMGvpS7PRybtLLjK0O03B
ObYNVYNi0z++NuHR5NSVQ5IXvLwMA1azTx9aNG1R5tC9jUFp9Cj2MM/7Hm775BITJousw9UZfJr3
uSCQ1Xeo5WCLPIu4wAoMVog0pr4DlBnDd+c+E6mrAOYYNa28RkJGAJup7FQmlWB5/FoePexJLucU
SS2A2F/8nLHFw9QyqGfSg5O4y36DNe+r0A7bDWsQuuPdbn++7lgkcRDe0hEoZwLpPoT2sD4QCbL8
JA7FINlEfb9v1A+4yspYCJO6pnEpjECFeubJ1+uJMVx8eCd52IlhMwNstrCcjyk1DWHNoi22uzG5
C6LdrT1HdJ6DOHIAqvKaa1EQ4UEvwGGsuIdFMhi+4hMNShLnK+ewq4qVqDggoKHWmxkm0yWPe7ip
Xo7vMRtbltMEuDYtv43S9+d/IWHqDfeYRQ4UtZr8txqGaCF7g2no2eblEyVyB87P9ODxostDuya5
Y8IJbaXYaKIYlapstObDUZc8i5dFSUxV1SRZinZwHTMhvuBD6NWS/ERZTBjsJ+BCFsSCghnR58Mm
BPhm4Ftp8ygKqB/6juTy1MyBAiS+8YExipJdtppC1owJZpecwJm+SCT7tXfOfJc2v00PRiHmVzbZ
oLlhonRhLc25hPmPL0z8w6xryBVdqk48YIMu7NkzmxOCMmaOBYRbkpyuDBSHDBwJ7HESGeeBcqSY
9A/WrzSDFOTxo4GcAn7t73VOviD1pcviV4pR+4axTaBWiCzmi9p9NkpPZ1KwE/otvlDMhB7yumdV
qA4MTLp+NuuZQ+2TNxFpi0GFa78OCI1jawO/3SneyBefxRfycr3VH/y9iKxKeCl6W7PPJVhf4Irw
2JfE+E30RjM19315d93minU1N8gnOxp7os+d4+3ZI+5cX40uZShhBRmCIHiCeI2mc/QLYtQrwuh6
calPSfeT7/DArHfv0evSHSzXhraFQpXav/pdojtRkEAMF5MaG3wq4MLVtxf0uqcTDDZsjpIfm6sD
E7GVQg9ttd50WU8SBe0mmE/7mmgKm1LYYXgsng5hQK1E9zwOGU8/tf8rqQJ+/KJrQI7rNRoUadIg
4bQgXeW4ZEkdZIpHDOac5PsTSVRtMiETvgJggJ/nsAqNwhX/+5ONFOfAksDtpOiLZUX2gw6a0nsO
9JzMlHz4MPWrhYjFGGaA27B6VSOGWTyPB6XdeaYhyHTWNXEIGRC+otctpm0WmfdLS7NlB5yY0Rhy
bY4Wi2cvbfbQrqqUrE+Lc65tySxGrwUtcS6GkEXoDP5dDHlo5LPdUEE70sG+7RQ7Zlhu6qQMfIWY
PT/ZKCM9sh4u5rlLGc0AN0+6oCVOJyZZ8353qe//JETXRgrocTbopj2OUi89iPqwl0SLNbiglT5A
gCH9IyOorF2CeZsWErR1GSd+Lx73X4fVXQ3eRgjYhzrfoIRtDQ8fW88NWgznYug/X+8ApqHKnc8T
tW/UPEsH5gEcXqhrnRMHPA/bbosWMTBymCpHIaBEJeiqq9YqJANGvQIRg4D/572SkCdWsrAakX2M
CkyvW16oUfBP4UQ7UFBReLBCmOCm9R4fAfVQXSMLNyHkU9PSL13DrIXLgYBasHgBQgDgAHQF2GSH
UvAaXuWqa7EB7klD1NRV7GLeCp6+te02Livt5p0FZNG/a5wTUXaWyhopZIS7LQBabS++K0oyF7gS
sd9gQ14e5L+9+ZrQq+AEQkHGjKPjcBctwjh4KY696uD0/7pdd2GWW7Gu1Khh8CQn9iTrA0mPYlem
qK7KkpNgabIALN0bS5rPCncdqvnX711mncgjkyKFyKjbBP1agYMxDHDyJdnQbphNcyE5Y+dTLRfk
RzbHnl/+q0dK5Pf5ucYrqHEZrhHn5BIuYY6Uq95383tesq26o6Fwc7e2dSJnMh2FNW/z6KBOxuTB
CRvcJJgbTtliGPoWp9FU6lR6RDk1ozmUhUD5Ow4LBIwyNI6s7l3g2icUz7TDiydgMiK+XwTFJqml
tMFtyJKSti/zw+Lgg8HTF7QyeWZ76L64exbb/NIUI66mLvVIo2Dl7fpVwl0Bk0Z0hsZnFX+VEA/P
zTslsc1y6zRUGy/Z1zETwL0oNt5BDYXI16rCVfBZu2BaVjcLSpoF6XoHzOBrZ+iM7J1D2PNxjBd9
5DxKmCHJi0NTeqbfp2t7S1ag6yhBxlk0gvUsc0vaa8kv2e87xsXsx70urdQWnPh6QlpEEBSqj4ot
lJZz1Tdm/DnlZqzftx4QNWL2//tgjHmKPCOrn2VVzn2NETvubPHG6sCUGL6KnFszJoLy6OUlXe1J
R/oi2PPo69L0Q7cuOy0fvNiVq7QqBrpalhFpHArmIDEI+eswkm32tRde57N8wezv6BB2SfgONyvg
Ph3ixQ4jySYGn+JZbvsULJbnPs6jIl6LEgxpBELilP6LPWGp4yIj9MP4XTQuxKTICmMIiVPje2QY
mkF7vRMNadRir2dvc0Ezb4q/FHyviSP13C6VatnqtOJgajLPt8MtEPjrJ+eSfogYwUwax5qYjLFH
WzTSKYvGOjRHukr8o/N10YQwjC4xVEHSuhnovLsjCPJFllkBkqnqeij8blkbNtujwNg8NH6+oVmK
bqShWavATo2+8v11CaJo3bCZFgfyDsb5NpXs11P6sVQ0XJnZKOyUM9A7ih5xW408G6RB+VYQoNXl
lxhsoP8mn+r8EDvW/5Bvs2zPaAAI7xk9rNY/szD16NfOUqhT8gl6buAFNEIxfpqAcZh1qwKddBz8
jYoU+tdy5aol5wG1+okiALE5ToJ1Wws/+dJHdEl3QurB0JhAw4imifnCCFaoccIhP0uvoCKtfWxH
lYezvDTXCp0h3RuyNXPWsAhTeQkXoGzKezkHRh0YRqvOFLno0ZMZWNUd2nQAsPUVI3htb6CIfGCU
MMCgSx/8b4JkWYbiZqg7CxRdYAqEWvqFJphB8aA3C+zu0sB7LaMBoWBbaYEGmBFGmoJvRNnaEGX0
jNV5tDQz9IWe0hxKly03UHFjpRhTFZacw04V7GDB6VusBP4k4JVxmAO2Rj53g2H7aqsiuHPL6uOk
Icw3c7UwbNMt5HAnjBgfgCISJm1lmTQDa/ou48j3ewS80ryRxYsf5cP+3DH9cyzyZ/itUabhS7E1
ETR3xU7opn0cIBcj60J9BsOk5nml3BpsrGbEKrU3M3lh2TSjORZWEfEXT0a+iBgRtdkBGonYYXrF
FYbIzoHc6VK35YZpqVALITGxzzexWMrkD0J9Ny6yOFm0u89Vdr61sj0jbB6bRcbDeKj3ypjgNgt4
flZ6GA7sgyME5lst7bPxKCDs88qeXYUnRoZmqi8PADd8LtLo7R9yx5rGEl4qRK3uUdWIeF2bUHZd
MMU+YPfFGnrXn83ofrJaPrDR8wAdVzEQWVI6BJVV60MmvHzBCAiGqvPlfe7OiisnJ1slV8kYwm4v
Je1NDCuFjO6ckRhOOJTvenf7ysCzSSXEA5qkSmoaOWtDKQKcxQoGqKVEUdVJprydOxHWW/K4Oal0
6/PEoQoTAPi0T0Bwi0/W71+jVlnBsh+X1iEvlBK5P0H7oo0p9/v/NGREDxe7BaVr+69ZHY/7XWSm
DvuyPxdAY7+bTuuOfDpJR9dZzhylD4kj4hz29FkxCvLZ9TkbbEbsrQDdXAIAEY1Qh0D89DX7VFN3
69xXM9GF8GZ5vCeh+wHF37wEMlorg1RDR/GNGaWoP2Jp6/lGedoFqRYYjv35doJWmyqGqJLDdT4H
9bq3newxmWMcJVU+OY6NDyTzizYSoI66VJu2h4/N03O+SL2w5CCo7ZeriUabxGeFKR5IXuHAHT0V
wyNQoeZ2rLhelSuA11U376q8szWwNhg5q1ExXSned7GXKnORjncOl7cYZ25DIv9L9/vmWBcLjAiL
m/9hFnlsvqmIxozKdu9MWhSm+z4Uc6ZFJ+Ydxrw2AnKtx28tzajfU9Ohl91vFxS7aE9B69GfOj62
oWlFFopxV2kyDnqzodg52zAcewxDVTx2YUk3/4798Tn16z9duPH5gT4iO892AxkZVZoUdJwbxcGv
Hwhl/DCt7UdsxArXEwMcQwTb2H5R1Ov5uyrVwYSBOgiS6ge5MuHLy0xzOgAML4aGfl+lUuzbJ/cv
7Bj5RupJCtXKoS9m0wwZu00iTKI9B3a1srL8b/9NdavZVOIg1FTUeOAn5Iek4HCW5bbpOddZCJeE
Js64S3gbuNCnzUubE/9bCLdljfsqKGRKtHW+q7Zmn/9JCik3QoyArACoAcZZyyuZXJkqoqAKQhdt
fc9p4fyppB0HzUbCvxk8jrfxopVyrx3SWnzPhDrVqS4vTw+RSfRdWroOvOMkC7KwY1ZKAKIlcCaJ
28n3uE6+lNolRTBl4Yt94qd7Zc8tX/WBbX6y048FseNWwhdw/gRiJbfUbF3kxU7RZERv8UHzjcrh
kedPC51uhn69GL+hUscG+lQFAnA3kByKBUpom7qr5ViPEA+dEJQdcfc3VfCCQKCHARaERM25RTks
yry1RSLpXXUBZ49gTmokL1kYs5o+tBUABr5A5xgKUmtZED90QvZlFg2SS+SZNy5aKM1dLdwuVyPV
ySNSddQFZ7/zhEDtw885cuJo2untOT0oQwdl23+Oz91NWw4KQclOYj4j9Qk9dpL1LJSlQa7xqIxo
qM8pO5n23B0F0YALu8nHrU+z767LtvCGlnjMhqxFyvNQkV8OgaWf3vvmc+ZCSilC5oLp98i+9wdj
DBaK6UU4s0ws9DeKvg3DnJ6qh4lXPCgZoJuweqdwPAFt96YyF5U4KOYkiHsnlICdKgQL7khaoFor
5u2McU/ma6UIfW6WlzQTC79pQnZHpZ4jP1gAr/p3JYgkxKuaTpIPyQK6IpLBTPworrlwDE0HWUjS
T1oPIPAko6mLwLZEsaSwpn/DLGOMICgjPofUDalt/4usd7dWbdsxPJGWm0M+IdaUlf+A36fncH0a
8U8Et490HlMih7Zuq/w0ssV1HvWf4Dvd4gb9QvZCkaDzEUTW5bec1hDu643ySGIk3B4WERVHvLNG
BHHv5vG+8p7YKkqfPBiSkzibjfKprgnu97GEjlGp6kXIFFWMClWKZP9xxbA74JeLzaj+z7iv0lEM
BMSTklYqJee0QkuH7vOVhl42khfMSx3x47f2PssjtYa0Aunz9DALXxPQ4jNmiCJ5B9iONFoNoAJv
ktGjrWvXKbcAmHzC41YXHLBrZqKp/aE4ZsG4Ep9BaTrFPpqcUXih2Mxrc4dclT53TSnS5eogYuD4
mGHcs5EnZ0sQS6nGBinRj5ZClw0sHtny2N71lPGB1mrW3bkqUoiUqnJw9noidPRKzIMQ/CTvgFqR
hPQV0LYYQth1ziljZui8fBXYDdyDOQNPZ9XO5eMQXWWX4bws32aOHQZ0K1Ge128bp9NQFPnTuVTy
Z9eoAC80XQIx2RNupkci7CPEfb6wY49KsPlhVoer3vn9RnZF4bU2Y1F/6+66zAWI239U8z86qgoV
GISDj4xiIC908vZ4xoZdVuB18lnVmkb8cvHVZLV3HgiBLcqF2eaZHUOl5mK/BP8qgDUKLPlyBqI2
jKvXQHKgD0RPGDnDx3W/kcrv8tiKACtzbLyyPoMA7gLfBm3ITE1unatVkgFxC2cDvejnESk1og4e
BNIW4DucmVKF1XTLJLAVk+H/rhqAwUXRHERw7EPNuHBHHpWW4js918KxcpXn37tFBA1rVaEkiDbM
ggbj3VPBKH+MZwYSLuNOXj2Sz45gd/x+7sxLl+vzGVNdEaHCdQ4UZsfK2KIMErSyg+Xb25sgtjLl
1kJXk5w6t2HJNBVhaaD0IZxn5MtLUTQKlDpwuQAhZaKxatw/xpkk7VZ2nT7poTxIqHkl+6Oeiu7X
0kkPVfm4M14rXYeigSimTdjHsnWWdbbEVN9VJOziHt7jawrC0o0yZqHRBPT5h3AhIrZHUvAeKM2F
kfIfQzJ2UZhezJ1oQxOM/82nR+dB/vG3cvBXlwATYhFZu/3d8vO2vEReGq0WIJ8lTdvL7pA47/bN
GcrfUCKPIL4MUimPR8IkZZKM6LbMT6VRTK/0gIyO6oTTxl0m5ImBq0OLbuClEc1h5xUhnqFSoDlx
delAPQ84AuCWvYGrunHEmEnMfnJZhvmdw0aG5i4C3DGc+hV4lzQ6T5tvOQgvFGTZo1fRbsCOeBfj
vO3xZNKun36kAyrB0k7pAY4HHx4dvGkJtU/te+FfDRosEuFZJ5Kcvvql48dtKmPCj0Mmh1q3F9Kg
O0TgLoDyVhwMWDhliNdIm/cy60LAH7zDzGWSghyReBVP9u9vVgMFkSDjkJ3V9l98pQYDeP1u420W
tQkVKvkdl9YOagqrgOl18EuSO7Zqk/dDHBPtj1gQeGpSf107Q+SKy/MpjbQ+ZJCSo/B0WAEGT9cU
5JNjr/qZIVoSAENjeQoP/aqvf6jtZ8JY2TGkBDFuEpxYpOboAJMNpWyL6Yy5PNiIs/q6bidk7ktQ
VEbnh/y4iIRUkKp4e9TkSTU9i4O1dTDQtfiHxhQqYt/y2I807QpNsB4vlm8gxRJmbP0nFkE+QULC
6UOcPm88KdLot2fVztshFtfxHnhUMuD27ggSER18Uylkk/r+thWxgCbKKXWavKFu6WT/zNUPQ/qZ
vGRU5rlK8KTnzE5ivC/Q5mh624pD2VOJCYEhqSsMS9k+0bUw0oAxTLntGjabui1oHfcXDcwdi88Z
NQylmViwuR3zDp/mJr4A7WXwckAEiGIDvGldrLgMvO4xrwI8lSp4vIARdTU2N9VuN3Ny5hdv4PeG
go04H08gG9I7xsQ+tp6Dv4DzN3TbG6TcntRZImVU/Zw4gUHq6gkK+v/oF3tg/qT9namZDLSoigW6
RXdpAYsk/RqysFmLpS6GeKWkMIQwCMYELTDTre1mjpesmrGELEiZqqh83tAy+9i6pzAaqyTZCsH3
vpqu0SgjVkdxfsBzHEovk+rF2DMMmfbNv/LRHiuwlcx8mNqoVQPQufoCp7Ni4TOBv755E1JCb0VM
xVb+OdYCPdc2op3xu9+B8W6ok1jQs6ew9y+vMZv2Po1uKh/3kpRpy5IDBJQ58WqkyQpMxvFEXlaB
jra+hergJkbVLYx5uAIhhj21P4Ndf2YJNVKXj2ur11phe7LDQXzbhq/jjFeq/tQTykzJIKDKjbnI
Q6Tej7PD2q68cV8D84G50jC70a4qDrZImniTVDa6RVNr6ul8AfdDvOCPlHhCPiSidyv86Lu8Myn3
Y0PYazzxAdvsIbjrJ1cKdDolwx1nKuImGdn8VGMc8RXPD0SoQKA9nf8zDXDupksUQBRLm3p3evcJ
6C/4q/sa67LHZNPgwIymSxLLx0cWIEg/5psz66p1aMcD0XpSCwoQfp2OuzZdqFgQhSgs4wv1s3dk
qoU/y4ouTkCUMRgYn0U0Klpq0EpMrYHyOlWABZtt6WAgneFbHjgKRsYjuTtSF1Axf+IzBQWYLkfA
3uy877+EZflnE3zrkEeAQMD56TzEwVbh5JTk3vEsOMiJZdyk3kGDQFYkIWHGo9HfaePszpP5mLUE
yFOBHT7qayHKrcFBK4CE1OQL7Znx2t9Wfv6xCap0kYiC3wJFJtv51+2Wyk/o1Ny4hL97XQb3DhR7
mdXe9dlREmVwRbyIlOf9zkJXdyz7MtV6OUASyn+GVX+hTpeilyeB87hSJB0g4vMfkEVlUylb49Ip
H+NDIHgTExfrIhapuAtUa7KC9LjHphm8YyBlFKdWIJ7qOuaJM+FIAWMlBVF8FlrlswZcvoUv/W6r
YFfgFUnJaSJ3vd22nOamJsuKYJCe0WlxTIiK7WQfjVQujiH/ghzZ2LWoLn44R/2UzlJWTXM934Z5
j2Cz/oU5o1NIsBzKC06lYSmSm47EsxRDmVwYpkX0wQYcKTYK2ck8b4xjktAd8b01bN0B6XU6VvWX
QWE4Io4nzQ/sTn2CDakaMOQbKvzSPfElzCRK+nSzXwaKgIAJrg+w7DH8t3PHA6M49gg1wPby3py2
aRvo4lOMiywKOCY+Jor18Igzl1F0tHoj1fZ912KUTBwBCZumJy+NLx1+ryU6sSMj32oGFfn7vtcQ
jTNq493nDEcYM1PV9WDIWd/Es/SS1bCkTVZ9po59NN5cDpa55Sz4bfvMrkQbacaeAY7kENU/2wJp
I2HV6n6gRP4/yp8tnPDN4vfUMMcQ2EbPlpwm4JSlcwrELaRtrovEn8BfNEaCqozAXxCzIr+MFFLx
7OJcZ/sTEhLvCIBIn2dNrtqj3dwjU1lHTkc4ECeClBd2dN9d6NeKZkmToVOYgRw4ZgUMl56F+RVF
XWbkjLKGj1lVE84zWwUgmwtwTpnsG5awEskw2BvEojc8a8v9sNO/ySRgqvdh9AepS+A9ymFL8HGQ
qMGaJOabBOLswVYgthnuUKahXtg2wErfndjiH4yCbjLGI3SpMykR+KWAtpge7OEK17zb7JmF12Qi
Jg78tUChS/tuPe0gul30xwY1cVxex462Cdw+q2D1UOsqhLH9wReIOQ2Gmnc79M4IJ3KFMWG7KAwY
bC4yGeyg934XBCGwDApbUyA2w9VFbGDqm5EPADrKN8cSyitHrMz5JN7XPVX/uT9DU+vtM3kPMEtb
Bp16oSmNL8Nik97+Rp3/IAo5QuUsOc96hbXU0P9HesHdsytAWJAHpDqAVameIiXDsZU/2R/ajMYC
Vx+YcUwHauEo3GtPHRfuubQxLJ4SYkvZOQziERwFzbVIixq/fAsDW1FE7U0VOL3kTn77jjdXjgAA
jeUTlUlpRnihU8Ls9c6WaSuhLXgRMIrOCdKvosM4fEaucNH+/s9C9CgQagtwbZMl0yulvSWHLKkp
m2PXUtiLiCvFTuqov/crfGvwfT8IksAhxG1XUfUlzITeTXZp9qbPeJ3xS+vWMyChAs7rQcQ9rZfr
o2P81ZWlSyoBklP4jqP0V6VtlUySD5qPv5dYl/PCBPwiRMNtTCREj2zar6alhYOHorb3BSKpsjkd
D8sauWkONaF1kNSnJ4y2HaWoP+tyQz3JfFTO9Ca5cdNdLt3QfKfCw6PUxvluPoeHnZYAwqt01aN2
Zyam+SyChzkR8Fy3xP7kRO0awCeNiPAZQ8xL2OVPpPWHkfWts6N4D+kTTzvgdTshba4MSyOaJR8k
a9gzo8RHWGDRqKKT+nrr3yXI+a6ETJLiYK/yxEkuRqRBamLmSPiDc+koKcsRtvwsmiPW0YlEUK2Z
kJ9dHp8bY7+IW3zwFWhieLVwvGfd9a/iLmppqvQfB6IPB8jEveqtJXx0u1Ud8442xV50QWvBXELz
5xPL4gZZEmU8sm5LvVQQnw1Beho8QxT0k2oeZgWOBjeO9TO+da4/sasCJxeSuN8h4TDL/X+i1WRF
NuoLzPhtoCVVCLmxzgTehWlEn0kKpka9KJVPEebNdhmWY7nUf0CHiUi2+tghrBI1kifmpW44KrF8
lKvE6q/jlEYl7vYU2bFV1SwnOKdjMR4h4QvoiDV4isskHSllIGcfKLyq0k40pQistafdSGGfLs5M
7yE+JpH668h016r4r8JlI29OhLhubGynF9wx4umCAYmN29T5s8TXHxooOvu02a7Y7ydp2g2uDG+I
JELCR14/TDLBFBItG9J97HU5YMEiO+T91cqqgEJaUxST7flazcAQqva2YNNECqwG/wexs4cAZq07
2of7+Iz6NSY6gzFpKaFswiFMpkIE5wyoMHZlfWCOfwMoMrVMgVG4C3o295iPawoN+7nDL+PqEBO3
OoJedulMvFCf+QUXz4IVdyTeh5ECnQqkwUqDHjDK0jUlShn01AShfiBC2KNcoJzpAAaI9u6TrFSZ
hEOIRk7BPFPJTdf8wT/Hv0ubqhMg8HlT+AjvigZnlbDmIeOt5uAXxugLw5ywLwtpWSRMHUe6L51l
z4EEfY7Jcs/y+QVi8v/q4Y3vBP9awFS+4naGGpp0Nbb5+XdWRIsQSQPad+s4z2c8HDkaTLiUMmhB
CcSZC/Rx9OLmFavqeHdldgO9sjq+8PI/NeFJXtKMINzgg8KiBQdzwWARlCifQLm0NALO/1LNUdvs
th1sldlrRqQ+6oCmxMwtl1u2K4VeIadYdMwqr1G3BIw17n2sGXagQINr9QbvSP9pykQSe4kvG6Ff
VXBeU+QOm/9uLQwMHZKB6etc/57zxf5J0kZC3IWLEBwfoiLGuAf/RrdOjwSFjHXX0lW+Im9yHAhw
rnHTX8A6E2+MMmqH54E0dHitU1LE7fbY/0D6wX8HgjT0ZXN1Ke/C8wpgcBQTQrETHlIZtu7SrCQ+
TS9UdoDBhHZknWvq6GFWulLIu0mhk531fVR5QhsX4osY3zIa/GrHWPFuO9CXN4c7MhFr8x42r0AP
LPYnMl0SqDPYx9vQh3qifw8kiSiQwdykBT8G/eN7uDgvpEaJYOlJASXWJimhH2UlqP2bynFDAr4O
gVZ7CPP9jOwlB+X8gWoxJxloPLoJxrdTtj2L8vn9oUX6AvzkvxJbPy7mLgCgN/eYnuImv0SEuadI
QXP6/nN9PEFw6ACKuRiJSbmtdZdSEWQ0impa9/mAbYCSDjqxgHOhxOW+xQLX8cAjum7EfDkvtnhh
PhbcCMTRkBRp0487/sfhmXG5EMc7VFPr68IBlL58G1m8z/xC3fCly+gyg9PfPsYnLpDQg+l2Io9f
uiPjVSackO7vvu8Yc4bFNkzDs8vqsQEAjH6JPNQdW3fb69E0K3bJ4zfBhBcoiifO6fx16cPiFg9D
774mwhqYH0oYJmTDx0+ARIkeujSFfjCrhk2Elgu1/d6lMuClDHsgsptER69PK0lKw0gHkVmsF82S
53ItNI1xnaHuoIq7Gtax2LTZaCK4FTDSv2WxApfzVbtX1feU143uErH4DiWN0TAYRlPAwlui9cMS
WUI0pxIzvSCxSH7NcxoiFAwUfYJbAPuaKigpUqyRPhJLxZ/+W4xibu91M86E/Y/zLmMtEIL54Bb9
E7UgzMB12Up8E5CvOf+ZeQjoFJ6qz9j5Hryhw5t4MwVyE3XtRPojv6NePTjYcolVXx8CTS2toZ8y
EzHSbqb4p6n+h6NkFc7QNYB9+Y9O6OWiB0F9n7o3z5YsY7oDoL/KYjaR6yltOUCPEiGazo/fsrJm
JHQRCXt/65x3q91KhpFiJlTDgEwhmC7bCCGjGBLneUyMRz98FZ2iwzfanR23bH2tCUKaI7QfKPJz
/42xLnDNp0u69I3T0LjLiGbDQKyI9IQ2hmjaxHEbbsMLT8SvUQwm1OFPImSXq9a/AYSNs5nP1ajd
ag+LWVX6h29W2CE0m+F2UmBuEFJCxmIyDjYASXLel6uG95p4O6zlSXbfgSFtuZvWVCobs0BRYSJQ
x9mLphKdXlyc0bNhhnJin6r608kgorlrQeJpDhHxwatWYHK4P1KadUV7MvL4emj45LVzKogRVGaZ
Ck2PlTYJkKXBZonW5bUW9LsrwIeuyTFzprgAZ7O4VUCaDoHwm11vFkPqatB1ngzPZOBp+OtFIUUc
an9zh35TACSXfqHdFBEx0fcNg34z1F+08fiiuWLs5MNxNysncgJLJlSiR49bj1ktC3iDd3wMwqJN
/hcM6omU1fSA8WRCq32lgX4I9lZ6+hUQT4MNixqldYUed0P0/B78rB+Vcf1y7a8CM6dsR4tjI2yO
a/IJvtjw8jSzpMEDuGyL4Y7t9hNq2Ivy6t1T3Hb3X8BfELfxkxXudOlCBPwvgNp2xYzFzfxyT901
9NYyDzZXq+GrLxVvrNGIrIWw5G8iEItxsTJPyLIcmloxQ4ToLRipML2/gbKw4Ipq0GRLIexQeHv8
f+z0NbDAgklGkDF3lcC7qzcD6NCBaL77/AFESz9FaLkZLQDq6CX+JepMa1YKuUZVpFD1WEt/FrEK
4Ouk7c1QLowkJYsA2pOFMn5yb5Kjg8xIR1Zv+oZjSoDx58M2E9zCNFsl0tAaDUDvdeibvLsHpO7B
JK4zyEon7kuK+gmQDdlnx+aiYjwvdcjzeyPZSIaTGeVh62+qINCAiKbXh1Utln7u4hTmyauE7OEh
Y5iyM6nDqDav2Z3WIAxOBPbbpHMj6iCsFVNTpdA/GRhP9mXKcztf+0EkFj0NCn/H2jmnunfK8K3J
CMWCaJHQyQp2BDrNoQ3ylWfY6WykecRkczHGzwgdoBsEMoUuCLQ347xHHVfdGrwqO0IQ61pIrTYE
5Q+cYfZUgHaB26lHsVu25FY8y848+LUDVQpn+55fvztKYqMjlKzYANZWrSexfqs5XBnm8W6TeXpa
7GcaDx1Tkp/0FuG+xhxYNW7U4BG3FKAlF/2/8fu8LTAq8Whkzgs9EpmO5Ci1JoDgD9WJ0HTsdj/V
9YSocALFSS/03l1y0Uj+r6UJ5a8nQXVYXaei2TpUYOAXyUA5tsj6CP/g3RX03mTwgTmWTmOd3YGy
fNL1mQHgbRSX9g8LtjSR0kzBPps0YJEMC0lcQ4O5/Q7yacqJIc6YhcYy0rewysUw06P/FWnmtdYA
82kEhTtInqp4qwt/Z5AADSr2Rum5zxHsyFYMqDkMnP/jE0fyvDbv1KbR8Xt96CrZv+r2g8pF/rPE
Ns7FzyXvNgLyAnMC3oU9P9PFPWgHjZt0/pV2uVhc2nviwIYeTSbHY3hd/vPjWF5mnNdCNbkfR96V
GB73yGhoXimsHzgB39Y/DsmH7Udz+MHf3PICmKX5dnhjsFIqIfnVD8IKmooCU/UlsvZo8LXCYfTE
js10tzQT/S727zGjGaWBzyTuU3jW+kpHwe2Om7OXpw/sQ20UV5OBJOPV3+/fyeVbHoDYmL+jX939
yHBcoy640e6apeYxLm9qYZUxMJGE9mxM0xhM2W3gVBciEc1mybh4ZaFs9qwEU3aJIjZEt0i68UMU
tA5yiISD3Jqk9qrP3p9+7Q5VMG/DcXimMwIK2wVv1CHHSzXlc9cWiV0zD+DhpZe/O2zwyYJsF+l7
zExG8gBzr9d0mpUX4IoCFV5m7Etw2CauHAPv8BCU2mT9oPgO0MgeCTb6RWUsoP3j+6HkVqkiVsti
Byf4KoaCbLJ3+rBdJ+198GbeaKWLQaIdDLFCEMNWGWgVeMyJCdR6nbaEpBJLR/kJN4IspUBmvGQO
iAPNHsosLrwbi7mur3CtMwomr+lNyXbapbxs9m5EFu0ACFTgY4GmpoB/aO8u3sZl772s0RUhRQEo
bMucTmPJUFxd4FEfUECteiFWWxJJg717TrBBs7YCpwvnH3WbbY8Ixbgqzt61m3D/UJKBohCu95fI
APrV+7Dn+Qf7Q6XkAFeZ1I1ea/7081dngQmUQh/oyjvJt49yFaRjI972oFCdt7I6QFvUUEDCBSGn
Oi2VqUd2pK4n/9TmFpmjP8Q2ZZT5RSJxZ+5ltZO6weXVliBL5OfZL0shUKVGxG+cOuB3qkvg4KeQ
vRaFYZSC1KbybzUxLuOdPgOLZaW2I6raJNdNa5RP4qBwYUDbRJ8sK0uHkoouyjU9Ytea/9NIVgWp
hSmMUlB79ioEGscZPwcdDJtEdJBIUtD9rkeNVxat2UK4Bch2lJNSSqdE29PvUfQR+HU/0eao7RXt
RWVDYfsABj3fzQnH2ehNFggAb4XN3f+JpxkmAB+uHIBDWRn+mZ0O1wBKh3FmRbJo8L3RqrcdRCi9
oby1p7DqgmBM2KRXVx58niwTJOY47zZKlRhSCo53pLBHTcZjxVzF6EW6m8BUUyi18GIF7IcFbnkX
4UAnWqc5/Z9iIO9cJ13nVi54a/1JivrvQgt4AElgpo0trYcplv8HreboNyd1/O1zaUocCfOsxOB+
smZSlRpPTExuFXoPvH13afPwEucMEuUUbK1hJEIa4Lf1MLxl0k6wFVXBT4T2+5dEFT4x+TThi/DX
pH2iZtnaNCkDCuihrCrMgbyJ2kQykFtORYXfJq/2pWNcu0blJe7wnFYbLOoOXmNAXfKIZAvmJBI7
0XOx+MDoIffvRS7wvB8yXg0AghtzD3mI8uOEukCw5kRvdvoRIQEYnKTlNSOexXCVTk9nAlTOO0Ja
dEcTIcdIjFMiBAzoDifdVBlVUqf/5gW9O8KMBuyKAgoIbb2/5+7U2xgCCuv1vaAhX5m8Lsnt0iTg
RcJk+mtOH1X+uOaNrtDnmGGJknV6TqbC5s2fJJv6cIHVocq7qcTCFy6TZcSvg2EIUyyIzzQS7fR4
T66WN7WqGmadQy7wSdZMPajrBVQ8PG0tOELl+yJvhiufNdpMIwh33eYvgFVr1YGBiUVputTDheSC
oEg+7CkayjpsRP4HdxY83Ml4LbFy0KPFGeB/u9oK1PS+9QIliV0qnpRPSSnKh1GJFzzXO1tHyr2X
SYa2upbROnVcb274djj4tq03vl3KyuQblBW2+8RPaSJqLcYGGfE7ok5wq1ozmyd0KPZMKPzKC5R1
D4hOxmghZhH8gf8+0a4pXxJTZGMe5eUxoYkP4RjLLF0NgUeU/M/jdvuLr78/M/uL9k7Z0DS/aVWc
PaZ6dc7pXZ0H2lhte7Pj8JommnBbf1LhJM2aIVRJChTvim8qV8MZJY9lNs8PpR537jzl689SFw0i
UuT+3cAAdmIGhnolr/kO56Gd0BPgn2O8lTtFvp29TX1iHejMbxB1Mam/9xtUCZ585C++RuBbkXEx
5y10w799zXBk4ZUp/Fb14nhjSDk+EhW78f5D1mTVQFzdcu3CW8Noq3JGai9VvS7PNDLgStl6jmr1
xthrzBZ7tQvyuBNqCu8AFwn2kI1//+mzhWdPKWrJ7jFkQnZ4+astGEQb9SIM+bl1eHthzxxfTIUO
oQyI+sKdc41JTqwGR04pPA/4TO0WeQCAfGJjun3bU04urWKMO/jFa75joHrTF/kHc1fC22mem0sv
xNb3cyNSwf7Zcf6nlKWMhSlGETpRfrB4xdy9iNgzDlPzickvSbcHkWj7xBuD7Y2jB2hFluk88aVp
vdyKGovXzVQnTdOYTpLfIH7r1m5e16e12I7Xt55N3pmEBzAbQx+Fyj3MuO0HGgvIuTfnLfU2l2jz
n7PnuoVLRBImenZ+e1zpp3TVbWBcGnMnSXsXFrhmk16dEmNwEU2St70haoYJ4QnNCBU5qGFB/MBq
KvgZ1LrPLR+M1PGV3rE2t/ewMGOQ4OcULLMZH2SlNFgaLAZLqz91ZH3wU8zFKkOpQUfdlHXjwSoV
EuisNF2uE+S11kkoa3ITNytPJpCOrfzq4UTn67vv6rTRiF4I5X2aDsTPV5oAV2EQS9wQw3gA0rUH
Ng6kDDH4eP6W6HXtIhMLPvstURqeWUfE3vNcoXpYWX4j6HUL17/GVXLTYQykNlUrorMtP47HPoE9
h9WyQfSIPLL2LZ8CCpjBfj+li0u17XbyBUt26XG/NWbMcmRIrlkt4+b7VTUH/Zr0V/r4wOlqy9QZ
4tRuTCBnjypHy3JMPBSCZwk3yfd2hP1EAfwuOsfA9AC5aaGhIfIpsxAgCW/skehLn0x+Qa0hRwDr
G3b+scvCuzK3opI9C00bfjLoU3cyfZbhmk6DyB8jjE75XNPJWxMvndtGC9ZCltI8qWApn6a4D4E9
aACiZvH/1KWDQ5ZGe3nh0kam5tiKE7gE0GMeSb0yvclirNyYr2rL9UUa/sTMfe36SXuKk5sna9Bu
UCD6M9S5OLtelzl+UIT9AXHzBpd0vje8UlKkgxG7FZPu9l4qDfsschaizoyqFuGGwsoAhG/TWYAR
I0kiR87WubkRRD8WpCgywiXMC67WEUOi9yDxGH3DxpL7qfWVWgBo6vOyE0m96gkaUaWilhDsoSno
D/WZCJy8UaIIkyd8E42i0mkfmYyT0SOYSKxw1O/e4ALceTvDpVEV12jVTsNRmWtL/vsDoLc2fLZY
zg2/d28TKXej/iiRxJw/nRHsZWIhFc4tPYn2l8D03k3HFpDHiR94TQC77mO9350lVI7T86B4CCuD
sr/ttdZvZBLixKkwh8Xm/p81qYfptq8toxRiCz0/eJlRknXQ+OK/ucxnCkHTkTd9MmO9Bxi/W0QB
uGB0HrMQpTOpgBPqVOS5DQFuQ6KH50irtECm5XfLX9knK3IuPtepq0Gts++DEftHrVQ2e+TR2nZL
ZsLHSSPp/7DZHJ2PApRAvrRQn40pr0VpFNRODh90pYsz2HW8nsX5mKOZ1489B2NXb2VfvlHzVed5
DJxG/oQo0rnyJ/fiuezmBr4OmlrUQM/2aHqyVak49wINK8fbVvbKvhK0nXsxHQIxJuIk5az9aVhy
29lqj6D2V6Ubyb3o5xmWS238k7v+HAj6l/Ov6hX4/IW9QNYYHsV9bQTCcszZ7XGppMd0jw6A7lgw
2cvhW9BT+HfMHsJCD8H+PWBRN2yvWO9cHZYaEq2uXymfJ+XPiNFLSqSI9LrvFjpJyC/r/GGp6yUx
FZxp86vzFHSuayyrfNP0Vo4IUJvOeitlVIUO3ue6Y5AmMefs/DXagkk83WrW8u3A+fULW6yOPaPa
3gg7Su3Cyg51U74dfXjnUkkn/yc4v6oNY/sBkkmNSzQeM+Cmk2elpd70VALpIOORgxvIRsoO7O+l
c1fp8M2Nmbl68j0bPRuoexl0qj3fed8ml+5pjFt1XMQe5MFzn9SHSeHJ74OzAesxw3lnHssZ04m/
Ci0H0OdegTtxqea8FKR0NN3UKRQOR3SbP0K+MhnAbjROD/VbOemzNpadT2H5PF2qnJpHhNlRoKEP
Y/WGKry+ibIBPuOEnelBbln7qDqjDl7GY+sptlSpgvgrxn3CfsEE4qbXcg4wCuNIvsmVDhmr6t02
FZdG7YQj5dj3CdQ7uGhhkUZqoHd+iQSV3JRav400ajulogj/H+RyUgQSy1GqGPzE8YM84P/IhDw8
ewc3Dd4xtSix4y5pTxG7TF+hnk2n2oBtw8ym9zTlD95Q+cdLQ+QdjYhRfFfhH/pVQhVSwOZanyga
hJv3iEyr49bdSopxqB7+eSq7J0Gbgzu2ypIjWLe0SZo953n4KubE4vAkU6dmTYfbVPRb/ad1BiRO
rcZyjnlMZJcckhmxIzxUcy+Y5m15VvsPJYwVnMqGL+YusPTODn7AvohumLwaVWU6x6cYUlLfwx7p
fQP7GYRx5UJPLx0jxn9PsowNN/h3p+JjVwlQvUmHKcTt/uhLOfTizQLrft/j6CdGBli1sT9VvR6j
CaK0SNvTWNBkGS4QmPGo5rTJFvC0/QsdLPLe0v3siZRk/X5soUYbfhjwef31sBRY8+QnrzU+BCJy
aHIpgKeiInDoXH7PXO/7hiAi5XiTbm2SvJXWy3BtGQ1zAluNXvRgBYe+JxMd1XinfuNlVgSb9Cln
AmNFHFbWbOogDoMjQF+0BuvakmGcPfQL9aJ4kFWnJTIGGhw8JPR1irk7k4pTWhkiblwWLAZLtkc8
4pbnjDGHVurUhnowkvo3KGhtceWrSUNK0VoG+stCuLP1MAOgIxIoGexjXBEtaKmpJEkBfFwYYXZa
zsJyTGxiwZ/CMaGugNJ7d9p7H13C11IOV+LwnR4tUHuGaDbIaEAjB2TAP5IySVjhG5JS2Em+NKVh
8KtIFuxeQQ2wv3S6bKS90jRcyBWf6g4gkNv28QVhPhGI8CqIIVQ7uCQu0aR8fwavRRFuNtldvT2r
rEl6Hr3OJMwMcn0NL1UFw8z7FPOYFAoxcJtX0JdLHqjXTlbP1dyMsXSJx/bM5F6bLMM4AklIHje5
FuVttFsVmnMXdKL69oK/+SOxw0eFxO6/IbN2DfnOI0/ozj5d7OsdhhuPN8hKnqA03UWKD6a7hUhT
Xr4x9xDCzbCdBLEt6kLWvu75z4eyfhhO9opl5FPJhtTl6u4nzAjZ2bBsLUKhZNfnIS0L/rTPZvWx
EG/bSWevTZjKptgJTCM0tkINWXsAvQS0jtQYfApV5v8tpL/QoSIX8F8EXB2xnVv7YurPT5DTqyFm
CXVbSxUDaxU7X6auCHW4ndngx2fIk/ZmHL8YEbktcSWaQ7ZiE+FR/1Xdg6Z5ebT9fQl6bccPrBC1
AH1AHLlCm95kXw63SrgSWr/lBSLPzD99TfKmMtq528DXM0TldznCPgmcR5epRlglhxICmdILfGMT
gZPsF0dvD4iPwuJgGYhBHi0SjN8whp+Yz7fNdwjCwRd35PD3Ayz8bUihW/Y7DQYdNIT1LpSJ3+04
OgcW6pnZ2sorfU/uWQlgiiSynyS5CLr+h2ccwe4gDBxjffWPCJTRIeTbouDd6o+wCfnnPG0i3X7C
/0Fg6+x6j7I4GRJGxWHF3BEB05ln+4B6qYL31nAEY7SkbUk7w1s/0P3vdCTXCkoPJ59zAocv6Z2t
9S7O1UVlgyUq1kZYBt3gEk6jf9NcTxblrDpeEWMlh+g0xnb6bcl2rSYsB2dAcG572CYtddSNpo4L
aY2BGzQpDDBJT7D9mPk3jxuxOcbbFsIXYUvC2s42A63HlO2+5d9p9p+eUr9NSVrOmR8g1yKP3RyP
1nYyAbWI1YtnIwL7HK9VUXpy8dUnulbt2m5lazBAWQXJzdgE1oydtY1s6Z6FhzgRcHPdomVxFdiq
EuPHqz0U6bptVUB100wWkCd7LZtVQiZvonP+aAAXx38J+yOPlEQu33FHoJN8V6KWxTg8cuslKWj4
C7eqzGJ2+H3LtKOHjXX9h7PoEg9N/bPmf+/OGxA/va2mXxExCDSQjEeAW/vyVoh2qOAyJHSeNku5
Bw2wVTVqZ2s2QgEW1PgYnP2K23VkoYWvPah853YOjr+Pl2Og+FKYehkgNhng9nphcVaNLtvgq0+J
bVmN3Gsa7t4UYCXREXp7Y2KX1UkZxb63R0I6j7EwpMV6v4wQqjqifm3g76XfnCoA22Z4s8VLHodg
Tf8oLLqJRGHo/7p811ihNrMDZcR3y00sa3c6kEnQcl80I4DG+9wNzhVrCjDYY07pSV0oe2j9k8mh
YPh2dLOa1UdHi0SgEPV94JILZfTt0fW5SpC3duOvCgI/JckG+PxV1iCiTvj+wLFr63fwLjwIVswc
7IlgrDAh1X/uIfo8jpkWMJWRAi3cJSzqYR27wd5G8khXIdaB+xeOJll3bP6PIohmrK8Mpxn+nH+D
AO98v+Em+kspzHYyIqR9hkHSwhC4j9HkXc+S3se4j2rmlJFPPBR/us/X1NxmQ9DfzTfMSixDmIUv
7KPjO90x6bPS5AZPOY4V16oiRE2dip6yppBaHzPHNN6o14GrCZrlS6NlWtR71x4XI+q05jF3oy3p
UObafmnJYL3yyd+kyXrqTlxVRufD5tAqC0smasr2285HsTRa0EeRwcsQPC8VpnX5wXdpwb6NyDz3
lSYIj+6SMlyewQj+Y1O5r5pBVdi73yG16xM0fR1PX22DphoEqGvp2DprwOpJnwc8drAjy+h9099v
isZzlP+ik+Wto9aBr12GAnFqFYmFloAuWi4DHA0Twgl5rj6OhNoq4CfBTX2KD+jo+JMewGE9ACGd
m32BAlNr5erbwWpu6Z/Kt8sg3ReYR5fN8I009+hIUpH0qh/r6xjDdkAQKlhrD8jkCYsPyEbzlGY7
cLs6/6n65zh/T2Vb1iTDvziK7BI9ApDWpZJSUhu3R75roVdPoBm0j5XBU9yIfI3cgJXlO7O7Auhn
GcMoR+NT7aD94bsEUDc1jbhFElZ3P1ZP6+yzMdUURTu0iw9wfxnUAI3bY3fj+RFM/okDa2EsGIAe
Hl+y6OsiNkXtxMkbh8jCpLvQbQIs4GcuF6cF/O5Fzx4fINq/mor+Nhyol0ZPNzWnTMlJErsi0Y+L
sI0ebHvttgdzv9BB6CjerBzZCpY2ZSzitL4sVtt0n1l5qVrP8HI5KsW9v0bSGGYJ9BDGTNsSuG73
k44wXi1hE721TExXnPsgwCL5RoD2eAW4EdrJvQ6EtrI94tV0MwcwTdxyQieiQFlrQYM+bpYHvWiC
E2YheidMmV3Bad+ub+aRcxlcxDsATUElz2yvgg4eeaXxSZ3Vo85OeVLVWCjeNCtp6Drj7VvmhbJO
hZ2RPybnxDMZe2K/vBfp9V3kTSNrqoQPsI/vDMLbhkudCau0hVYW0vxA+AjPwOai4/awHDIH2kgl
pHw8kiswHM8CMJ7SeoqDZ7id9MXbjKVPFfB1Ve0sWrlFXdd4Td5q02EubdYO72yEqANOJJoJrzAL
OdeU0wpTm5PgWJwGDJzI4+DHHmPBe6diCpsmvO1vzJ8Dc9EXwOZLY3TdeKfWeaf/Fx5aXXKDe5+n
43EDPdeOnxoc7gFAZuOZUi7iMBCEi5ioV1Be0rtWlXdVmanOIW0+kH5SJOaaM+e+LtkmG5m1TWaD
xL9xyHr+C1nP8rp3v6r45d1Dfklv+BWkDezylRn8+KnHXpsNyDDLhrSwS2CwloFdmd1OlUIKwrd0
ZfYO8HWuMAsJWmSy4Pc8MGN++YFAh1ekaTW51YSo0C07kTK4YhnFJp5lUKWhQmUlfHxim4uIXRrO
kqe0JfTqMx6K/ahhSiisAWUEMY7f+Y5kJk6Yfp89+kC+Kh3u03Vda0AHtksFxrV0HKe6kCGB438V
Uu/q5PDQ1GmW1VSk+G0N7bMBdmIE8W4kzwGSnMgWR5RRHhraw2FbINhEo2HSX6Y2EqjO6A4YDcGI
zOuVjoXr+xYMOThvoXVhFSpjrCHW+U9tSDiDeuTLsfDFCtnBK02FVpcyOQb/YpWfnzWgmG0n6LKx
PXrAL0uJtdz0i/MYhaLEC/XVxyZD5D0wj4btWZ/r7JB5GddFX03rUq9sjvTZTowVnMviGm1dOfE7
akfnFN6OcYDjh8/hq8ipwsIp6DDvUFv3DbJuFcgcc3kD6JktEI3bRmxFYBIThFyOL7UqZHCr9mZT
7wb6DGg+XLjyjbKDLmRcVRtVczZj0seOlTgsN7dbmv+j/ltB2r9ur/jGyDEZKmle++zQr25OwykV
Tcpc6bnn3qn0gSInUTP+7ZC+JWUIjdKFDODn54irU9VcULSeu3cAOWP43iv8riaxlxXRULhi8EsD
Mxl+qkFaqe05I7NTfPpiWQ9UEcJZwaUqPW+IOL3Ub5o60UlxCrYqHBpjNvNsR1qh8ke8F9uq/7nc
CqDhaOJRGABGjjDJnVBaAmWkTqqa3iTohuCWlUbKy/AqJ7BHCrecfxJ2tCqyPAc5XGFOp+FwIg2h
xqQjsx/Yj9n8tu/JdPd8XMQ6nhEW6IxMh32FThGWUBjQ8odb7q8t50Iwp0XvGBosboQnySiwnIcR
AcvbaHOu7SxVzETUcK1cx56xow3/seWZnmQjYlvIxZKmA6EE9kprqC9xfsiLjruc5yK/VEH7zX3K
2bqPp0MQa8oRFbzVsJKCVIw4FVzu4pzIXIrtjlT9QjuXnBFqpmRdPFA6xvWt8KHdo1oLLWyqlw/Z
1By+wr05murs21QmrXHv/Mx72yghOoec8Qakogh+rjMXMevsnv/AysJu5EA61p2iteXFypQZfB9V
64yMqPg0EfmAOYkFRAst8btG92wUoCHMG2yTW9ElGOTxC5JUwZTD+IA3CIjX0peyY3F+2I+HTlDs
aNO52YT2Z596h8iivC8dLhiNidDbK3ze6cWB41jm9W0CauARJ4504L+X0es4IUGLy+7yDnseNs1s
UWCqrZkMIHNOmMdfS4hu+I1TcHtdbzULH3tc8e7o1uWTOSOUbJwBLqHF1Dr93NQyly+dADaM6xOp
RatrYv7yf3thGATSlPzOa/jCXTjRuFY2cqSVnn1TnWLsqxUEMj5MKcpp7PvbBifJeXfyXWvFQ6x5
K2cAgZb9RqtJhV/7Ae59kDcVQYHhnxRTal5to2i8Z6nAcd+nhDNK7U4FUVDOrXbJ6MMhAAWxjxm5
/eMTy7Tswle+o2e9HoirPBrQXPimZdcl4ISfyVNjujyG6KzIcZJgBFn7ZljXIpaTTpMFFVgNy+BB
b+PbgYogUrGHX/2r6UzMfNE73iasGgy3yl3qmmfD/YKKlzmMvxByBVURFS4OQ9szC0gcp/A+tXi3
SN2ptZ0i3yQ16kCmOb4UTYQm6Dbz3q1yJFxDeGgoIJJ/9FAGBViYxGnVeTCexnTNeq4O9C+KyrmF
NdHQhh3klcIGS9HWJJtdThlPai4diLl2W3ktnl3cnYB+o8il6kRgJq5A1+XWXpAHNB33dg+S38b9
Vs4mZ/qTIhGZiRLrX9fwyL9fYf3PuIcPZhjePcCLRF05EFtKyjXe8+EfQgU3FEHHxhku62TpXmzH
w0YCR8fHrBwnnpy6GzmQgG3huolMlqwo7VcH/nwmgLF5XgiLU3U58z1XGfn5kXDFS1V0B0Zy87zA
aGDBSla4KuB9Cl7MTEbKX0gYPmjGOgSOBiqtwJEzYse/Xc/Z25wqvODGZ+NjUjJWDjtDHvocESsg
3vjovOEUB3og4xhmdszoaU17AIDowf5vlbHcmR8jSQjipHlzAJjL6rUQrPo/6tAez0zRZPvu6lez
lFP+Ead1QJi2r1XHfG3KjO6Dxa51lxlFDzvXZwN7ew8GEkRRLSlUdvyHjwNgqgZm8qzRmLY2yHMo
yybv4UcWbar7ZUPioPCNe6cAF9z9zCN/EosK9aH3lAMKrSaIwCTEac5jnlZ6g9mylJVo7YVuYxKE
28OAoHqGqRgXP7L01RvIDk+UFOipR8VSCFUHINuUOCljqeteff7EpANZCanrX+4MSjFmhdhlN6WN
nVhYngJYnjf/hl7PNIwV+8kuOdQYAoG9kSRZjXfbC3DQwpp3+sMZY+/S5XQRvU49Vu6OsQcb6UjP
4SfmORSF2O9clfDIHVynTk1ODwQfVq+JohrNaJStw+vmd1rVCLtH+pqVUsHkew6fjJqzQ0jKdby8
9eZA2Y171EBs18kH2NeBpIxi2SmWVXqXZWh9yvLYWQEmUioMvyIh9WMKWfGHGda9RmAh2EvzWQxM
j/f3DKxUQGUmA6ni/xI326CZrPAnbJSQ3OPxfMuwL1nUfhD77x+U26v4OueKHxCtvuDgk83hcT8I
NTk8sy+8OQQ7NzNKQOmK9gcSAg03zhHiM+wkErDqgFI3PzAHsy61OsfUtcwkrunJvx9cSUxDMXRV
HXcm+WwXPxXnIWUoGbcK8MS+a0Yd8UCVDilNlinr4XyRzeOL92E9OxcW5BdofLl/+HPqlbpR4xZH
7q4bPOaUPLvch8lgLWNmwJRGcBdAIhjdWAjPSYL4ogy0Eobqh7NEH2VUeOhb7TB6rCdnbHIDD2fD
/8TmLSXfhVSi7eeACHtDVHWVEaKJfsBVKPSaP3tFc5Uwyc9y5mY4sNOxHSAOyBY8tYnhsBwkH5zs
m5AJk6bRrhCxTv/rRGogVYw+RER+fVPf/OhdKAuQDKN1b2LJkQZg+lno1dU80PZp8EXkaJ/VLkhX
L50a/KMW3jpPvBKKnIpcxVt+CzOZWso044MkCZl9PM0fXl3wC3JyF/CqFhJ6XNTMGhK5lI3mUry4
/iCbzVSUQjl9hW1eC/8gZGc0faqZIPjUJw97zhlhFqZxmwpR6kL8CyhppUFw5ghmC+w7AFBYLqsf
CElSseMPC3H4vDD1rvOHJPK2l5/Jw6P92DsqQxYwjWnp/BsLfJpwGqze48e7roYdABAw/AccElv+
AibLtzToyI/c3cTITDhlUGsRr8jokXphvvZHLMTRB9+zktzWk9fhY8k56AwzoT7DNQC64NXqEuHS
3NAjK/JGZZ96Dy++yLUabp7AJJ8yR27OhIFf5Jn0Z2jh+iBGxKOzdGxaiHuh7Db9z2amwAxov2p7
rgQW0eiw+rvC7ZM3RbgbzQY/HGRVGjR5HAy525AUnB/RLGMGunxH8u8aMVfQyp1cVph6O/Em1rzn
vaOEjTXw4J9w/suAHOq9jU3E/pGi+bm8j61ymUp1nSnwtRHu5erFCwDJ/GMFhDpUpnXI+eJUghfD
xYs673WPmdnAViuFP38u9IyaCNrTh0MEXqfOexb7vlpMVxDkaIGeBkdIPrj6JPNRGEbIra8pSPCo
bBUruLKCql6HCN+PRO5Ia0pb97DV2Ky6S4rkmRZ6KLM+Ob3zMACp8vud925mZjJT8eBQ9tsIlRKc
IZPQQLHI2V6he3rlFtN8j9rMY8Rr99Dt2On0EMz5WxOtt75WyLyQRAj+qtJZbWs5N1E0Rsz8v+/8
xwW6Q4psokOklRXiW0SiggwDaLJEiIaMB3/YuAmkfP0csNGNtm7N1hXsvLRMtXRLs7AztArxfBja
4PALZA/q7PYrCSdsxxnRM7y7UzY6dzmDoN9H9coR/QKJ+Y5YaPE826Plh4iRSQ+652EmmFbC4d0K
7B+nDEXlMNeBCshu7AJqIHbK2VM7WSZUmmEZbtojPw5RIYo7qfVibHByeiylnBvFgTFQznXi9Kq4
rd9o7RFcR27i7t78LB336L76+KfuTumwPmvtGWx52Todqyegv7ex+FkpvXBeUNmR9483Lfix8FRW
Y5d4kvlGqoICqgHc+Q+gqY0TxAgJu+ikU8US9dzv6WD7GeMvVaIHOrzsh+erqKYvpizsnCb7xjOP
an41QxbdISwLuZ8Q2ELBBYX8AlF9OUbavYTEQ8GYp9Ongc+lu+7sty6iNGzYhs6mI2Ix6asNi8u0
rLIHyV1ji1L+N0nmaksDgbTGTJ9jVVIG9C7/SCLTDKGhUg+MupuUIcL8xYL8youua2/ttXpUzv3t
BwSTxKog+iPwZMGmMblCFZwAoE5fodZPiwpaLHkSFk3h2qxI7FSmZ9xCGC/15lLRNOE/3UfYwZUe
iClO7ZpZ1tf1RYlCy70+l4QaAwqLA+HEcoKb93xCHNXxvNTqnO7AS9TcPcfsz3j6Su3fCu2yQsEw
/5S3QLLy9ZVsFIE3timsMMeDSNCBQHj2EHRkVSZn+ly1oe57GMWkNBqtmfVxfmtddGmoVrJwGM4R
eujZr1bGr7V6l4/TZ6vRdLrc6TaJ4Ykb4Cn0yMbVFD46Qug2uILLex4OvdlvNm/+23+NS9TY+lvV
Rqxba+gXoOo4ZzHnwupnBGXraAq1yXd4Fqms4I1ZOY39lghvF2XHEh4k07bucawvTOU9dDvakJ2f
Sn1422z4DJAKOhYOqTDLgtwXwr/vhGDdCKjUkIFjSVhoyfekANmGtcSUqLTtwUJIu1UepGIN3+sm
1Qw0Cr+F7oTi2qLKjX6SUZB1IIqrdagzak3b4wLzzhEVeoZQSF+P1qyh6X8xJJTbQ2i/6Y/VFp4r
0q+CgPWv0sGk2zKC4iBS146iUSSmW2nG9MJcQ8RgC7XReYap2xskJNCMcE6xKwDOp79bZF7wPok6
r9yauv99nZb6SUnmmjOn25Llw77XdFW+IXExvpPkZAdsJenB5fHyeiIc65CaZoNNg8YAJPyo+0K5
VdEfHxZes3yJmgHwwzJEN6G8prGcB4ecHVmvw3vITkevA+BjjqjdDlKaZnhuKelHbZTINFavQtWt
jpDNOxu/lZcC/xuodCNpLKGc+0kuWPrOg/di1rIFhZtNCyBZvm397bZ/35LgVqrh/hK0vv+d5e4p
PF0FG3PL6cKAhrF/e7mR4NAVkraZtqMCvVoNFXuYlBxjfjFbAo8IPujpNILY211M0orSGhgL6L/s
v0VJeNA2wxKdvPPjJ4mjKG7lIAmlLWVwfx0T7FB+1IgDRFN5dCXxGy9jUxVvn1zoGhVxnmYh3EDC
NVAFp03g00G5Z0A5Iy6Al//fgZYiHYRY4z9wsWJcG1WzxJXUoj2hqmO3CZR7oOPwx+BH9IjrnagA
Vy+pPiyuX8Bbw00iti8HbYBfrOStoj39XOXfvSUii83gF3j5DlX5VU7n6HaGhwO53JfBm4pOnklq
RBoYY/4QH+gkG9vK15M7OdmVYe7KZEgfA1SteiDx+VLWoBhmKCKROf6KjSheiYMSAEMq2zSro9rr
2SmYxUuruP5j7YLPsi98GNHB+Isj5IZf6zKaVVUwFN86NUqO81LJuZvdWYYGUSeE36mFQ6VX/UT+
MHfcII4i2H4dswqw4fppfMzfBMuAaTMvqbPLqOM8qTiMjY8enwr5JKgPcqm+YrA7eIDXp+Cf+vTd
drt/L2nvrQZmh1iCplXiPEWqGsF5caQ8kSiaAwct3h6+QhPQTUtNJ0vhMLrHF979QeVumVzi4KHK
AbOv2/uqLXMBc6bjMlVDsMHslXvvl4xucUuospYTrI+aRaVNP7kPnuW3219jV+aB6EeedK4JV5+m
s2PMJBP9cWjIJtBBIqU7TKW9Lma2VPyQ0ZYyBL9Aoai+WUBu1mp7ZEPnnOu99+/t/yF95Ho87q31
xUngIbDJTXnosXeIV1DMVG9xx+ltXvM4CFH2qHCiB6P8hShS9AuSXN+3FcELOBJUMfIbbe4sWBVZ
Tu5hf29hacR1g+nxj17k4OtQIqe6O0uXvy7s5278HQQJ81t4L1H3G0N8+wCebNlscsInlWu79p+e
h+XcQXJHTu7D3hE+g9oBCJncIGEko+7ygqOAcwUsDTCPrS7/stpV8bTMbvASy+Xl7EhMXgSCKdk6
DOsOA9rpV7f2nJ4Oqe3tQM5wqZrP8vNp5gnpOgE4NST+3P9OeOCPlR87Aqtha+kcQAji1ri9IhNW
EKdTu1xKLKeLNzsqjFBGh53Sh9BXY8B9CPcbVTMYwWuUMHspYI+zGJxwFO8mXTVn4bE8KAK0s8Kr
258bmcRxY6khb266GAEy4qqg1TCXYzOM8PW5RWKIb9UTzP//QcVhrnXu1UMGdc7+Jd1rBprff+VV
FtmXz0R+CNxXy1uC3gTgUGm/zrB2WBoQETeRYnYBQRETEFjkiMhIUWlWx3aQKX+3Fc9NPajHmTpJ
Xcm8AKG1ZMRSVYGhPkbLZyuQajQlEVYw04RiIL6ZohQltcviQ3gj2bNjgt3fPCvZyqAMxyQE0LLT
rsYIN00Hncrt2XxMHGXZyEqj2CHRZvw0+mGeTAP4VNgWjExALqzvTSFdir9upyx8FzpWo7TbsSl1
qmPHhSkYYCxUGqCG9RixPFYHA/vkcU9+TY8r7qssc6ZFHjD1nqLqVyZex10esURpir6rwEPwaDds
rdWvys3t5zCp8JisJ5NLmGuk2r5kPPNzpXtj1WHped23ec79m/Tc4neA1Z3EaHg9tpOsVB/0Qnf+
DRvdl+ynCORk7ZVYDJ4FO+NMbATp7q9CFR1ux+TSQpqK4y6COUKFcaFai+cRp9Sp9iHs6FsSKx/E
Lz3EdYT2YIAbLhrpHdmKtT9oD+ffC6+dsc3n5sSIP0CpKeYLd2bUO2k6EMxxXXp2GSKtihtBIP9A
PkgxkRPxWa2ywWa/0DMVZRIeXohSN/nQtVsT9lHHHGblSD9r/8A6VGeKpzlJPAlm2hSnhDCZZTLB
UjPTT6rxbPllVIlOoB8OFWN02QSkWaHU9U1TzkfZ4dbXaQiiJ1bXDqQbH6K3IYIv5DFsFNGe1/Q6
+deTfs9LHSJiNOofUctdxjxrT9ek917JY9JTttAOFC22EJTRPYyyTB9GE7N4vl5ga3P/FvcTwFOd
jy3HUdn9L3iIg0FMjDHEeNu1ffWuu1PsLluZ2B/PNAVoSj9AsLsdzXoAigqiFwdtjD7iCW/4xGgg
eVAzLywVzoU11iK9/9F9t58/BYiVNHIkIfce9tZ/kXllkslI5/VRSLdP8qiao3zou6YzWaQzawBq
6sEoRG39LSzYjoq1Das22WnuyIp7A91tHkmftNkZwfA/MRtktgeG3nqTjzVMRoTiDts+T5A8S2PQ
VLZs64NIXb+xwF8OztCg3eSBggHxSJFChTgKvrtPdqt0PLMj6tHGGD3+R6HlNy9PvLNcMDmhfIyd
5Ol1eyxpFDyR07vAiNV+CJsUtOEZjJfLmPq0GDqj7RgWTvDRSWz1H9M+4dJpEHVVUhJA3U5oUhjv
lyzZYnIdJEeFR4eH4bXYYCa0PYAfVgUC6XK8y3YPO1CTiiPHQzlgJWp1pgPfdnQ3T5oZGtJEYyE5
q3YXn3I14Entz4GIZThnoYMpf8qpBWBpRRBpAH1/kQnWuKRgBDpyQcWF91n/k3p8+hMgTGTtNjRd
OD04yWa04d/Gnmh85909iLDCDcWJgTivApWPL16ongD9zsrrn9+rBsF14ispYm3dsRbnuevjJPSB
2O6zcczbMnVmj+6JXDbGxIye1i10f5cKqIjRswQdivJjq1wm0n3t4NqThaH6WxO9u9zJ0jHmR1ml
9uilAc8HgCJ6s7hVcGsIDWM0mxWLSYWASVlVOT4ZiU6MXULKFifGeI+ZR2UlRjoz5S6p9whmvcYP
QrNNBQ/bgbuvF8mZM1+6NPxloZvtz3BdLdqi0k7mMTvAtJVtLrnvidz9uSvqtP8a6N0A+tM0hDsS
5k0E5/q1eLTqf9EWHtU0t7g13gb1qI3vG4t/A3aR+31rA2K8PDj7i2CIEt+2VfTLycr6Yn2hW3EK
d6myXgeLR8s47J2VllSXhMBYmzWjg0DXoITa9b1o/WQJf3hcyKFsuGowTqzKdpD/JzKnF3jm3FJy
Bkg3xd65d+Q4gMS4B17/aPBjslTXfPpXpoou7h1XrU9n5lZ4fcIm4Zelc6BxyWYjw0hUlNbuJ8Yj
+eTc6l9K1IaT7BaRuGBjdyAxQM9/LAAWKD8DQcxTNvroLl7zfJB7Q9uAudN59NxDUc42yNbTdKkB
EDtW6yOr/poCkJWMhNiNVWeBEcCPk7+0l7+FAusi8xLZxdDSQS1gV6hC1uldSVw8rclQLDRCk7AB
ipNr2eBS5i+/A2Fdmynrcur1fAtvGtyOKGIEEQJxYGiohb6fptDbn5uiToJATGCVHGdwHejmO9Tj
XRQgosClgrYG1bsa+QGFG0KG3IwAt99avU6lLYPry7NYcJHM2ZQNmRWXmgxGHFLhpxyyVeL0lvjV
63G0KWOKYNImbPy1RDmDis8rbDCxOScWI+hh01AaRMhXiLw666zoPwbAXD8WM1iFeXpDFbcrsYTp
JJV49LgQ5GIRHUPw+LhwtCRXGx+CB8n1cHutz3MfKFo854tLXjlJpVLWS6Y2pobvYJ6ivKH/P9AN
aNr55qlFeeE5sraJ7v+s+9AZM6HcaRQ8E5Ultsz1p+isrKId5t/BY3m3l48b32W8sGe6ppRei/zU
R9CDIaYmDzAu/TB/HNzWN1kUGOHFinGomj5amZOojFrbBtSurZS7XwFfdVQcLDYYG7zXpYaH/Ccg
xC7BQWMwFrrv7Wa18TMew61kEuAFcCkoneAFd/Eco1m8qVkXyNntWFMgFj53HBLQsaRyxqnjq82O
AlpC3q3/GyFdd1JdBx3HjxjzCYl7zzft0+kCH4ur8tBp8Nl5H/dHlK9BZGG/XrnXnuerkCvLvG/F
VhmhUBWUZix3Z8AoXwCgxDSRlwzdmDCeDYst8PxJWnhgmZHone53PuWe0F/0BcXeJNy+DyiryPJ3
cvygmxmHmR0e6ntdk1J57CPiWs2WU1Aznk5MUGzF5J93KkGiNcaCbEsPuRQQykmGcVvCumgZi1lT
yNaWPjmpFmG9edXW1pF3RSIRUcJmD6vKnpLVbERexKHlmTBxBvSB6sNr34Pshx4cl3LuSbqT6jRL
Fr1x0g4DGqj241KKJ1dnkVjRGqaJUerMlFDY9IALu8f+v1hsIat1fSs3BFcODUA42trrElS74MUh
0KXjpFU7n6+byyuTVBzmwkO9YtoVpPoDYjdDu8/qAc3rlnEgBr70RCrYlN5JxGpi0eZbdqAR/nu2
jMZsLssp6+vzVMDCDCYa5caMPbok0KDUTkGv4cYULHltFpS5hxLk4bXnZZdcHA+Q3Q8LK9ApbxNl
3xTlRgr88WoGWkYW6ZWSG/nKDy/hAl2a1VVnjjTxzYrjIHKoVySu7byYuhbgE/vtFUlu+LRB34Dv
F1HtSVcsf3znVBeouBfvB4DGhK6NPaSuXipkn0QdT0Zl41JuBDP2psvchKga3fACvVGHHLaq64C+
UDVMTN1CH/I6jHm/8Y1OymSUu0GD4oTQC5ebMf3etruTOQoVR7S4ZOmNF9fWvZuto8Vg9yWT3fz1
jMrjVfu/dwWnu3+jWjV341N5SOQ4DefgJSx07KPeqz9bLSvZFmsDYkq5p1ADqWgBhvfjai1XJyXA
5k6HfUYfNGhopTh78jDi+qP3aq609GPkYYAvh0tUA6pLGfF8m8BpVyp1QVPyWyyZySbSFqUsxL5m
LF31Qo5Jc2mF4QsVkO248HPp3wZqMxB8wgaZMQgOulMajQFGE8tv7BSYLPvb6wmsM+sqIKdInAp1
BGuqr7rsOSsojZboZbK7vmz+pL5tYT97NSm5W/ZZH4Xa7feFP3LUEXenwI0s14ZY4y5Rhtlkwk3v
qmEh1vVqnKcveZR0gyiN28F2KjUMwOgLzTGU+Vbv5Suu+MSbOQ7QV6mXGJw0O2dwL3T0GpFfOdDy
B4dcyzZMAs2V68DeWHxArQgp4FtRq1StRYFHbeQhbzI2AfqciKOzB82FDO6tQ0PpMGAcouKYeXhR
rvTza/Hotca3GPY89+Vu0Y0UuoYZ+7afH4hv7L8arjP/Mu6eRnQxqwXnE0Fw11nh+1gsD4lCctMD
YCJ/2LEW6p68GOF9/5wOGkuSyrtJnUe+vfWzpq+1t7PYeh4ZnybxrwGB9GNd/e81+vX1gAKj73Wr
QF9zoz9SK2YdpMZz0bqH8bmMo+hTx4HjAfOgP+CyhgscMjiQKfPAgKs5SHlNoLHRJc97DQnGTA4Y
LZJK2VXsTAKYOo9Mci5czNJKsKUCK9tFOmsfhhI2xUmbhuCl2aGgNMdYaHLpUxh+jxJfaB8TdVt8
LRgzeiw7ErZO+HwPPF3mOSx615O7Dh5tX91YM92b8jxuRcaRPYH2tiAA8PXmm5xGbQj3r5RyOT4J
7gHsAHO1YhcBAmMNxWKvERoH5zH4zKNAbZpubEKn8Qq3hAdk7MsAzkiD7HeeZ6KDZcV3pe8XlFoT
kxVow52UXhrlm/byiBCrpbR4LTZuU2TfXo5xbOjEctIzqADu7gz/csWPlC/A4tvmVUGcdpxshajY
9s4nGVnBmgNKgS+2vz1BLf2qzrUa9dV/UIeHfnJjiclj3RTIqkG7TzvHu0jj0okNB6jgaVN6nr6u
7CRRtJlrNAhaujYtoH/wip/LvpT9TnsqApNu9z1LUhObZSbQZl2HXVg3fE+hhf+vbE2YQSHe8zyx
Pef8J1uDb111HXlEKgjDy3WApB9nCocWIDo+Dg7GSbU2fupxOwu4SI8sNA+4K2fkNiakddDTTPh7
nxQgDNm3mbs2BycswaSRszmRan8/sIMYumWg5IN4OISZDSbb58cLbWzVM49f4DWkvQ0dW0/Jxj1h
63E6gEi39zKcCcOKfe4BF+gZC5dkvwid/W3LxuGBiZAuESP8lj0CZYnp9PKoxm62quots1r/SmZf
GiQsU5jfMf9+dREpmg3ibHuQQixUshcFolWrd2Z6g8fMynSySpildGCCrCoYFGknjTI4q3iB7xwT
FsiwdDd9QDa1DIePiBWWqHJDrRGvNO1rBC6ZEhdUh+SXo1CNzwtufGZAvowxli7ww+m2+BJwL5BL
syAznNrjHKtG6CCG7HfSqb+aarxadhbkOGgpeZ5jbH16ZBwbC0pIw6x6cF6k61t0ZeFj1INw/gSS
/dg17KGRUvfYyMKVil1CeC0X/QcNYcEaY78ruwfP1mk34auZWwvO2oSsJWI9zKYIJHRGA7ewy1fH
bxNqOKBbsHkjRjUCby5ka94nTAGy+4Q20VuXnlK+lTe1HvUahmb2+ltWALt9xznR4mraIB/QP7Mu
s/yH1D+avh7RnsWBOjfWvw73Te4nAdTHawqTGQ6Vjn1JcLmh/j5T16ar5AEbHYN9i+qmGFVc+aJ9
bDmC8Xo/zgkVicAQaVTT3fntX7PWdA+KiV0cRe3l0s2DqmLEgt9PtMPPpZl5ynUmFTuAvyo3UqcA
hb8n4PILHAsCyhme3VLN5PHHUH94yJbRci9BsV+GQ7g7s0DRccBqgco6h99j+27zOnLRbww5sCTo
kLBHBSFhNz8RuEO8yYTpRfw3ol1V5IFqH9gAPqJcuIIvEmw+hB378xrfHMTENeAennliTCsv8UPF
OJL/toTNpXp7HZVqdrx6XDnhPQueX8yZp2UHN54bXaG7E6QM8dNjzG+AKR8zXatGzt4boJqVUgJc
OwJGc5pL22QiC1PklHPjCBQlJXmu/x5NEEnA3D2LWsTHRDthWevgZ8qdHllW2emspAe7bJjQiZz5
nVRCJ1p+BHrrHH94se4zkT8lGyrOTDOHPn0o4eQ90B7wcUfhF2Xn3l1e02n4VQwGI2rvybQfhLds
/YRYnf3hbR0t8T+CFk/MzgizIg6TXLZvw5YYs3d/gnMQOQaGB+8MBBtqekmZzVikH6VICUW3h75z
/mMyK0K8zXALhcxEpdb5NjraodH4Qnp+WfK9HprxvwT8y7Oo1d+OJIl4xsHZDA9qIDqwKvWmkAX1
6nklh8OteIYo0YS2YajNmwA8TMMfMkc0geZjWDKrLq9yqqJ5crU9XnI4Ub/j9HqpKZutjd9a06X2
DbviQABnRDELRIZvClBk7d+1y1EpWPW5tM0+Remib3gQwe6Umqsr6cy9/6dJpyjV3zTVCFKQoRVo
C0ORZojFf8TIuH0EN1zntvo9EsdfjgZ9kbZ1oxDLi29CWXsbrsNFkKtZVpKckrJzMa83XXJR91m2
VXUaPzBQhypulA7exX5BZMl6Xr6U2JKXl06ZRVBWR/r+l51Sw5J0IlYi/08Rl8fQZWkSHdcaTaGu
5baidbAFM9Kn2ElKryFIMWXdFI3ZrFAtKGR8CnOEC7UU96sfQjWPW4nLS26D1Aq3+HMGPTWLBZcV
DNPMu0Zu0HHhJ9OTc0A4sgEtAQ3ugrKGLgRFaS2FHBr4wJVfvfRAgfofQk7cumpuWy6NcHZEYhtn
nL9a9PG3F/qTACA7hWPtavq0Cvv0jeFX+pbxPPPO0m5/HG2YPVLFXmlJqh+XSJSaE08HVcF4zQys
KZ77JdFgGI1jc1tW+I+52nULp1DqA5XQPqTgXnHObFH0FTdhTgLUKk8ZfpelxtghIiAIBUEkgqQe
Mtkb11F3sNMb/jpZ0jYAnaGwFKGoZokw+Y/geqBdjK9Ge5thXt3PSBMXtrVR9dchzrniRGBQapud
1iw9IzWCIvE1+5mp4O+rzBWCYAhtpNr0JiE4a6G+M1ufmL4Q5rDYgVpA6NeUdQM74gFMFfyZ2038
hBdHKqQML1Y54UABk/wxmgFWeNluswmtGs4lX8zPHTfJx1snzVqn/EHBefj9l+6LbE4rJBig64NN
xMTVg0J3T4FS6fQaY2fU2FpWMXIlwkcRqwWTpxGDdP/5bsqG910kXLBa2AYtAWsdOLBY3RfqIeGZ
07SK09nIuhZsNd7nO93hwrQXu9lxB5P30qWITc8yB4S+KxuktGCils38qS9JLwNQRvwwGKYEssmy
zdFruJKyNug0T7BsL/i4lHsTdJdCQnX7ZJpo29yFjYhSrN77nf0NyPsna3UYuBOQVodY+PPn/6AZ
EPTAbD45McHEchRavtXU3ezhDvvcEf3rOtditXsiUPFdJRE854lZJohaLuTcjA91QTarrT28jDxz
0ii4za8K1glBviLuoZl7BGkXA9ymnqxkUU60BrPFCR24RThPpuEKXNMWlKfcgToj9cShdD3ZusLd
IYYEVIDYjYFPE53fM334RKVi8nxkvwld7gcSmcdBk8Ki2UH00DpFd+HCQeuvDwFFeOPLLlBXJ0DC
xoXPSA5gpvJxvQeN5j0zTYHHLMt/ILCvLa820m4VEf1EQ3QdEJ0XSiO5Pz8vMn1QswAF44wdoiMS
bkpgTCewHRd3tJNQYuUzARZlQUoOhKTS8IliYmuc6Y2b5zrSGH3hKLKgNSQfLaAqA0q4/kIybYJS
lCujuPXCEMO9iCuNWtG9lmyBB1TrzbL2ihZpI4K7XmBkMeS1aX804lz0w4pFoPhrmpLqqSxzHiKy
KaRnHsqaym/v7gYobdCCclZdgctokBXaU/wl2qRTEUPEZL0cfKMXD7667Ov8nztMKEY82Hx96RRL
4AQYK7BHZFgwWDxTeMFe22bJFIkbjARt0oL420//7TnBrSxaFAeByW28JgjgvnXyTUxMqjqLRTKB
UNiX/Tj8AKpuHt1jee5pxm8eCRGUGhw5EF0ahliw9MKmJqs+zln3h0/jVls6CmkgT2ScNjsAFNE6
Z1nWYI2fAjKSwHH+hV896wEao9pxYrKozoCe/8s68jY9WSyyrQLgYBCZMtKgrmZkxEQ1Kg+3F6pt
1OXSfqi3K29oTO7g5amrCumb789BTJwYhysZbY8Kif5v8ChVzrF5QYZB3UKk8JwArCRAmSbjU0OO
Aun1ByrwHX+etZkYRCoO/xlfbwcjJo27TDrF+UpYvB0A0BNyqE/j1AyAz/9By6OcmdP6wV+nCtH3
bSU8OmAl+GGx9HdYpH2iu2nFxlfRGOntsraZ+VlUZstmpnPnUuSKlXndvrLfmB5XLW/UDRIO1E18
X5Vk9YhW1fjsXXx7r57fxFjzq2sh2E23j3aTHv4LTzDwqAipL9hUiRnFAz7y72oVAHhwnFcJec7o
NDU8GFCwhoQbok1AE/UvbGE4mynCqzFP/ExiQQL3z/wdPpLZ09LMw/qhCTxqhv1iazN9sMCdUtpO
OjzuUm60v4q4iibR2GoR4Ysztt5UqGGTDKhwdtAZpa4apFDdoJPC2xF3C+DWNUgAq7f6Br1dWvAR
qA+vt6QTOdVXxdfRbRPH8cA74ja+tuJzlvceoSvUsu5mTxMZbhPOYrwQ42cVq7zmWcyJVAONiivP
Ld4yBZt+LDnFqRSDDD485e7CPrvcGeoh7EVb48HO5fPOoCDMx+iGNWmojD0SAyomlMYK858pqUAH
pOr4tmGic7QhszWLWiip2Y42Cp5RC03rRVRNt4yxfy1irnjpg16nl55XcB5awRrFnDasmFIHawDe
rbZ2D++vFjmJhPY0i1YTqMzEDDoA6bJQ1NQutYVgMQglK5XIUWYx51pMPgt2icSfEmeJD3Hh91fa
NC4+3KExF5UJUPVQcEZW69YC1Pmny0ZaJrEM0Xl+2PMQMn8rKypXXYEaZJZqRyrcBodtNiCqWltp
yaytym3iR+BVddaPmgWhieY4/VA18utJ6H/fQ1iYJCSxF+x0Q8hin2yeCfQ9//Nqk+C3Zou6Q+1X
XrTYDTGY5yGAF6s0dKpao4A/imiTRTnDm482HqGkkdBOHRh/SrMKRQTBJoyTgU++5RYkod/BgKjW
ElReLVZI0JjtvydRoUnTAZuAb91bEYHmJSmkhuGC3T5tObClTvyNC2DCs74YVgHnpaMu5vhWVTb0
nxd/rRvOxyxULb+b3RB5eNKYWGSrnXNMOgxQoa12mv6oaPLUWCbk6UuLhezKm2Ev7l8QNAD8W0bL
cS9Yu5ksHoe0gD7aptGTDCWCL41AK1QV7ahk3q19vroJAob0JenK2D+D/da4UCbrWJHXUmU86s74
bIajjGTUxHLtoxKkeCLKRVNmRQOWm7wu78sAmVdmVBQI3zZAzuQGNviTc7gnVAkqAYg0FBSRt0xa
L/WT1LB3hU4e+YSt914RWwewNhiZ3hxCsbv/5/vuexFb8Tn+/5u8i4cz3CK6SndJghiu2tTq9fgg
oArKzg9vBrxgfUgK/OCYjkzjS1u+i3MUBZysIoT3GruhA4n1VVKor8xoPsvFkknFFQAXgJFY8P5P
FutPEyVNbBfnAbhxiZMevvgrHbYZB20UUZw5HHEDlLHKAKaGkXvnKAdHJzKMbh00geH6OqP0szab
DwaDA4wIT1wt++LCRriAowu7vsRJ67UsHl4JzblnJ82lZIDIv2mtdDHDj5IoHeA6LyQLZpk2hHLj
RQ48WVYneJFtXBFuW+xevoF1j32zUqqFXKD1j8w2qD2MwNwo8WqjNGYYqyAmRISO3oeNl2/Jpdol
GvSmmzyvN6B0B7fVGWovmnidiRt6Aez61JiZOSICnLKWAymJbieKDsb1KzslUq+IHjmxGGJX8j5w
58aF/E5E8qj00dExF6VAFUUKJO23wSUx/n1FEnQGQdO8TS8dRNrD7XSeNqvoUNxembz2Tplgswhq
Jim2HizMt3mbnQNLZS7Slr40gVoLE9VyhR/czn9tZ+9Kt5w8Geghg9/WZbZhqyeD2MGH95/VrMkW
Ug2epvPA5iB8QLEpJ8iuKQg3USjtwqIpi5LXrj0JMl1+N9rfhk/uYPHfrV/jrMRF9f8VAANQWG0J
31yp9tVdtaHDNpSDy6lkaof7EdPUOHYLVZ2030yx+1hrg6tp/3+RyXlbwrH+8zakJ2GP4ir/EHHw
6g+DJWJdBtfwy97F13/TPYAswH7FfMtER7BOl+iInmauRKXxSTg1FnLKOwcEpuujrnH3ygNcZULp
dPOey75Bgi6+77DABbZhuC4OzNG2up9vAkZb1OAixnQcDW9v14OF+FZIt5du6acjvyEUfXp1Tw6B
Zo+glezM68v/WQBaE9JkzsFp+vFI4jYRItCTMoKfTt6HnjyaW5vFP/FoDyzxpwgR/+DkckXfMTHK
wy7nBjn5bOqQC+aJNiqGpR4yBfV2u0nE4kek6CUNWM2RoJ99IXL3ncRqMqhDPuyxF72iqrRfCSZd
lF+cxNKImoeuQVDQ3cfg2xEM/6FsEasKUnXcp8bSVkWxXUtBsetAsHrucpF6MsOxS7ECslC4gz4M
10+uFuL0zWBtanW6yOLPJM/33KV8PPkbiPAarh6DSCrXU6Bysa1hoNyNCCX4E4hnqeik9PDdHtR/
BK1aZcjNzAeJ9LiDkooa2FD4kMEZSn663fF0MLdd4QUMv4AaFVlklKyNTeEMtmNAeblI39y2pR6x
RgnLQLWDmCnWZeoCPYucr/Ce2gPG9igX9QH9ikAmNL1fPnKtWRYqzUCQhPIYl/0KWKs2RTepnGiv
xZ+yfyUb0St7chbMkq5DnDtA9mkKcPx9mtB9AOfox+lu76BHc11dgKuUe/ge78b/bIUK2xtTpFd7
3B06uvjW3wBcRXLLwvm9p0LUmB9D94KsF1Hf4oSctXuZd6l3/WB09jGrEBHKOswaA+WMtCoxObiY
gU25NKeXePFGCSDmV6C24tl8PQhg3r3EuTQr6s3TPH25toeuSD0l/Vd/tpp2g4gXSfszHxY6vhxT
35CatBlyciipCz1Jz0PeIhG+eAIqN9gQNWQIrfwBlje0AjKbhb7u5vdoAernGgXXxB4/d0A/bqIQ
DxjrHfvO7Pa4BXIJy6hDXMfyttqu45yf2LH1J9RMzAJDmwNAA9EKmxRWV2KWbHzoOc24g7blDVYx
ayr9MaxKNIZzfGsqvoEVHp0EUJDKHVYCLfap1M4zkG6uqypE0t+amHqqTIKeiUZQ4L7rGofgZuEk
UztkWC4bYfkrgRY7Mk/KysjfUSC5HE9Wvu+oW8WlJjDJHcW6xxc+xzFA5rFcRzTGdoXUM1ljxWbH
Jq/ATy5dVqQmyH3RLfnUHQDH8lBvfybxtDkgSzsXNyayCZro3dvM/EYQ45mEMSKz6XRBAvigziAv
XWqhECKcrZQl2NzaloSt0AxYOLJQzCPMu+FKjtdEjrSq9lmfEB9rSop6zX/gslud9myiYYwNUpuH
jQH+B1Bo5rBxneoX6CTl7ILUMpcGOxpSD6gQmDezjaJJI0NZswI1ly7eGNH5vXhRBeUWAJV8JKcc
2+nLvd5jt0Nw7ro5v56tH41PKCl1CQnpZNq2601bIotU1ClWnuGuv6CCTnTdidMySORcBeUKnY2P
DLz3gvZcsqCHkH9R+9EAOZ95wBjJKHDy6YjFxzNt7klxHUXxfjrJhyS5PsE/A4xCvoKJtDbeIdki
7JFDOyl3BO/7NF7x9tasEX98kdNveYr9MDflm62U27CUVa1L8WcX3k+oVA1+mDXstzUdvICVfqqw
Aj630zihsZO9rQCCZYocNJzlQaxSerxNg2Fp4e9vLkfFa7zpffnYSgN7cAuYEP4Ar00joJ2jkjTp
matpErSCEqNb/6Fh8X6GZ42LZAP7SZf2i/2xGL4BGZ/IQ9HwPCQWHGimT9OnZSM3Ye6X9ueeXHbX
kKoAs/NAIpmrWZk3tw6jkUH2tWzwVnKqG3n/qnJeuPCaV1NtkkUJPCVj1VsAOKLeifLw8DNLDrXF
01x/koMQnTM+j3u1OWuyhX9XVkPaADrUwBlWS7lHE84JKjVdCjUFvc5LbL/N/iQlnLgcoKEjcEJ0
5p6t16UefMWDf35SBM+VKzBD96E6zNRPJ2hwqlN77G3SCKPuNVNaBxqVSdO5EdKnJhWmSX/+ITWN
kMvTEKcd+/MusrKUXrpdNsxt6AbPMKQFWgpktrl3+K4uQTdiapbQns+/LcOS3i4STWWu+Y8D4gIe
FeCwCIDD8rRwTQuEVhpFdEVVeUR+8fSj8L4HnH5KVlcBiOETa0AJWeK7snHUmWsyfpr0/veF4n+e
l8oT0OqAqkNyTpfqFFauze2Zo9MlBAUrUwmErWVz5t5wbAzJY1fcYwDhsWElR/U17+qhZhp5F3rh
73IateV08D27kh84l2IWmhNZnIRWyIl63WY58zG5veiwITA6DdoFspHkE9jr9enk3YQBtotTpGlb
n6AIvVKfINicBuqXeB0KVvyp0ElLU90K/XSdd8UpYVrTRoHHke7mbjIDz07O3rMN+XgeBrwo1xeW
P9m0szHKGVjoDreIKo60hqItqqT7I7t8SMP6SVkaVMpNenwTeVQpOKoE7sbNhA2xsjfKEG5g13M7
TW7gC+ujs4HqsNec3EpQV2QAuI82qt7leSo4cHxKl+XnT2KQ+Uo9j1X0maWCA0rKw0uCmtBlEx32
wLOzORyMzMIckDo3m/VDW4r9uD2SaFN4hW3RQq/1o3l+NCAmoPgxmPAdyyLCZioqch+sD+cfZ2M0
6jOPy1ESUe6vupldfoxF/p/piDN05BpFIyNSPiwN2tz0Dzk0J2IwwKfDJrxdu0TJylAelTi67Sw4
CWVnSb0UZT2gBbOic/sqpQoMTuGsMO3yfJe7lJKBZ64BI9EU5z5+iVP9YIOhK04EtqCt3DyC4hmD
OZ4UE/r7UtB+mE5I/TW2Fk7agzNXogppuyizB8serd57J0J8h09O2oFlMjzLvxiGpqqElmDJW7q/
J2ulvV6H2nauCFhJyt3wOaLSaS9W/cw+4AlBurf8zKrfmqrOZX6PHAi42WMM0ywm1O0NxCH8HBJL
ALwk4Ylk+enOpR/QTNr97uHofYgsqbH9PHRKTAkzRUgHPWoLBnTnTPCbEC4CJrB+6lgahcWpxVB1
6YOvqSLSYvi+zU+jpmbotple5+6BkEbKD4uUH2gXliyE7iYhiSC4ezy+ivfob+SkgzcqcblHTGTE
S7L+asRJURLeQeswWUrtB+LwjTFDpAr9zTxMIYcnjVKX+dT118rmRtm/SFuEszdWLxSEbPJQMa3C
0LErPHRqNiWnzqOQvFUFXm5NkOtcapULKhpCDzCZvIBG3c99J7g+X/PgrXfvqr+ijDVLrVb+h2A0
9cE0MyN63h2CRRHimBTanC2wIp2QOQxslYvAat+Tgfo/4WjIUZ1gQszXrixWH+90LobbI0wtU3Ms
wW6HWe+VR3K13TbyRVs0Qu3/N2CeR2/GfSja6r2YU44tqFBk7/iWegSQT6ogHjbUzl2naXk3M35a
mWEXfIkBegTgXVusgDPwNquGk7St3CME0eaHMDi7utjc9yATJ7wP6Em4ew28VorFj3vNB5eIs2ya
1vGCF8Z4BHZsNwqK+JhbIIns4afgETtFtxSqm5y3fK2M9m5WzGfWnJRouaABZoNCZPqE60Rch3kX
N5SVJS52QB6DOBwMVdwqEwQ3fs+EUHiRqyRqYIiu0klgG3qWBpZyHC+4k8TK7VX/lSC/dvVIafUE
y1l4u/tYncqKiAxouBJ3H49a7WBY/IYQrBp7iQiSVWhU44KplbHAVaAuF6RELTABzXlFg2/usTAD
ZrK0YOoQTFvc0UNEQ5HgQ1cwc1mX1FBLIomzFqkaOOrRkYwsAyr9IZvoUJ3AO1zDLWjUqnu84NCW
U9ECJ04vqpLeVHSO2/KGd9kR6pRZJRc1eV+JciZ6wxyij2+y1kiPw1wp5UPOJrgFVstL7qoaZlPa
f9VMmkR9qQvDCJ9JgYBQoIc0wZurOrrt41oxE1OqUkEbDof7DYR2PYxBz4OZEzAV24qW5yrD5vKm
UBwT/GWy16ZqEWL2/iFEFBFiEbZsAxqUUnhHyTbowDPs6S2S4Z/HUtN/gtWsRWCkZ5efB9wLI2DD
1qPtknQm9WkqvQXitDNVOrGvbWedyh2XsNtyEyLHCzuhyO2e2ApS4E1XKv2DsdFpCzpk/KXzuPYN
GZmH6AV+2sm1WBjV87KM6Y/IjyPMud2YtxTN+R+4zrTNmDBGCChqAuR8Nw9/LlNK/N49GvTllOwl
aKIZ3wL1scNJftlko5zaRFgnSGc7PH7TiAdvek/Beq6gMAPp49o62LHlHK+DV0EaZAi3pW3e04S5
08i8YsnygMDCZFF+Oel/A2v8nvcbje4RTTRE9nlsCONZ1xvMew0DobTnquDUV8sirzO0mMlbq16q
lNXUmQJVYiLG6NHMhGSZYdRP4hEcBxGnDPS7u5FeXOOE5+soIGfleZ0LllfIeSFS5pGa8udJb8Xq
t5PYtQChJ4Wt/s2gYUjQ0i5U8M+Rlv9e7PLRoG5+zeT73rrdrBq6XmxpVi7nwCuj6RpeBeT7awzT
HKNC1Z/d7SmmkcQAYFyDASwu2PUSEe4PHAvtMuwjJ86jvzwFXUsCdcZVaBCtHg7/ABfIFw8mNK5a
1zhf2P6nN4s3BiKu6itfCQLhyYZdxHtNuYVfTVaOqtZm/ZEQ2x52quX+cwN+iwPqh6M2pckjBbJK
uDPMJjpOYxwjznVTv4ano46i0vgsNqKuejHxQySaYjeOEjZIKoOXG5++nptDnONUin5eqbAu8ipM
yJE5/s6yuMkUKbvU+HSBsy/HkSSJ+briwEw/lC0iNGrhj9tTtv3i1XD6xaapRgoPmswqz0RlLS59
7OE4RpswpvV7iNjLZEbDzlWNTsGa5NPrTSPNEp+40M4i1JywiLKLrAGhkkLwNhcNxdtA4s5EA9FW
qvZfoGZWlBm8er44f78s1Vct/Ccs8AF+BDE8vKaj1zLFLVkW+H1ajJDfE+Sn9pv6cUbiNwnZM6wd
82DwQ13DVTnrliiesOtZK2TZoob51RMrlp786pT1wmjY6cpCaBV0oVBotDcRHXG7D27oOTfmSP/p
BNA+DKjqdI5U6lA1Wf4n1dWGZzwLPdnPZSPoaLRPIKcMsyq91wF848L9SB33p4EoUIZ2ZMWhL2ay
+AYLtqOPWLfauoRSqPXfOA6HQnYpWsXaHk923jeWJnDfEv3QRs/CvO+42YJ7NsyZ5tNTgjgzPXbv
Sw0VXQxbec/jC3svz+eOJrCCEl5uO7hg5bnTcNGR5Tq5v6A9d8OKgv5y8G1p12pdzvXeFildMrgf
FjBI/Lb1Bmnv3qTG49K99gKwyLNCdk/6VJAebz52LMjQDAJwrvVr9TprMepbsghY0XiRjL4bbx9Z
ePCgT/Pl5MU+25gdeHH9GAuLkCJ1/mrG5ijCETz/CG5SmtKo/dr+PZlil7o7iZAL4zEVbdth6gTm
taf3vkB7t4aPKM87VKDoHzV+RkXqi6zC7ojc1OSii0ir+svrt2iWhhIVsYqQArvbQGnSx0zeBIE7
JACzIlyQ8m3IbW8bnMZ9wLOenvQeY3qpeDMv57zCx1iJC/Xl43AHs1Eyjl0m6tMQGOU7gtoIfL16
Dpd6AG5F9DB5nWjEYWCfA4fF5l9PYSmp+5YkuuTDM3KJ9+37fF/yPjwHnsqkBAI37Tri5T7frVOw
IYAmP0sb1/XFYuoWQFmn5PKOhV3hIeLQCex+LcRXUWf4WjdQn76s6YgVSGsbMiMqnYgqd6RIMM9A
wmadrk05cctmi/LkmY7WO1Z0vJ0YoFqJC2Vcio+KoJvF1lIJWFq4HboNRSBXietMp/oewQe8k1sz
n0O8dZq82pQIBjFLvCSjy80U3+QtBOv8bhRsyTjMjMYwsAkjm+qokt5JSnIHQn2ymUlPb57yh+Bf
knldgo2q0Kh28HUVz8QXdJJf+avGpoGnBzP4joepMfuLYhJqfCvDLAhTDJ6axpdu3zS9cLayZLw1
Zj6GGTN6LBFoR5mIvU7P8y6tkFrkuGYzlF/3Sn/guKISWvfv4Ls/ec8CdIzthZE428fzb75PwKhN
oWop/5E5h3nbKW4gdX1fp4Cx/0HwpyceeTP7HMx0nLlgW2KHBcQlnAk4S40RihNqZho6pA8WyeWu
xQfYeNmbFkPw8z/XStjDRNPk9PXWzLN3V8JEYKVMMSGrX1sjixXE2iA0D+l3QD/x7i3c31VyAH2z
u3xduwtdVlEGMlbOufkoWHwzC/4MpcQZZeaVlVqMud8ekeWRRoqnEUj91ICzXpCkwZu0PXc3Wt/1
tFdWUAQ7lY04kU5dVVbcuJO9HFTriCFEgOWMZgeq/tc7ZWAaGTp7Kk4182cM/hXNc/OMR5Eq74fh
+6U8a5xYANbZBIzn/Y5q8IUX6a//tB0o2/OfgFviCvB76Gj+OmauQsTvXDIRebj2r33bqHUlw3Qg
o5JwwM9pEm50ZKaAwDslXYDqhQUpFTIrUnNooHi8xGyLuvjcaa4W2eG9QLCojIYInoqcToBi7RUQ
jKx1oobsm6n6JVbS9zkK7XgHxEfhW/AydCdBCszaZZBjpyouMIq4IMyoBNGSk2LqpY9E9NuBF9EQ
T47nvs/ZQq0zPPHsoPCuaJJtTn+4FnuDITEog9PBJdBCZgDKFjgTxtgoTnlkul47aguizhhwRYcp
eFCrhD0Z+OEIPfAgDFbLYlIOr/zhXTeSAY8IeK0RgPL2JHWiN5TTWfSL8TcrtWI3OZIQja3jwvWR
lSKcA6ZM+WLnbmMmcJMWxdG/fY/BgWhhjLyscQLWfbW7GGfFqPbf1ABIkdcnj/20oKaiBQ/907Qb
eyLIlmZePf9DDsLIhezOACmxlUJxZxbGlxyk++4atBW2CpxHwh/CZ1FHx2RaQEU9JrbF4SSoGjeq
ovDogJk2QK2IdfZtXWqK7fzgBrU2heAnnldO0nyP5En0qVASolHOxui0Avkp0NJDriHRzgE1kIUi
jRFMGgIYNpREijvbnbSxjqEz2U8PctHWAtd3jg5EZEL39SLd5PRqcACMyxXG6wemoyrba15iPp6U
TbIszaZybgvc1OHg0s2RO596y6dkWseDBQDIHras3AIgbfzPSbAmCaWU+dR71P9+r8e+6iSfVJKO
q66OewjLb/7bXQbnNxwzrTd/zdy6xK7jTGWby+AcwupGz7ums29iCKHp75Rrpah4MlPRq5C/IN1W
1DZjYHxYYXKUJNDxhmm5ocjC32GC9fsJUKp2iqTZi2EZ2So0KThprIMCBa3uvTJBs3+8X0MXf9He
n5/wIKxr9iOqUWGs2ZUTvh+TNN/QlULyM1S5AQZl0SczCyzUPlv5ivsZ7t7APGgNwOQf98BYRyFe
dRr4g7eq0VfBHNJQLD/hnfy4GKinUWkdHH8NIAp8CoAEb04RC+QG7nxo+8V8QYL+agp0Nvh8Ha8X
3NE7u+ALI3umFgYiAV5a/p8yW3Ti+jgfeLSd8oSvYdq9BBo5PFu7F0kEbJHyuOCzENHXFD3xfRtI
WrI4EWjZg4AeTohrIq4MnaJ/PAPuY2ZDQKrXia0pLFgfFLY6H+XIQ8LiTm6oKqzGkLZPbw2ov3JY
CZJ+lLTGwYbjrEgL/37y70CQ1ASZaUX5Ause7Dc+uTok2uA4tPtThGX+LJHLySNsiUfoCUdHKs01
r0oCINZXB+thzEGKZpJQvB5VleFgymSuu2TKvnvl05i/41a9xFrQrnMiNyv4SChvZoB984FgmjkA
OYzIBfNrzw6rSk32NENyxStG/SUG2JLw2WMynrgrjXA6cmyPQjMDExMawWTvqa+as7pr+xgSV+cU
zPQ3sh1bM3R75sa19107fpemzJTZunroyPdEY1DUptntnAGkPBhX04vBBcubdgjlo2nWVlO1Kkfy
5cgo6BzbMJRwIf7jtl+3EE3DB3ZIgHVjVLZef/dbcDvWqLTwVeezHg30CmZwoxE6kbP86OITWJYi
pnpUT0zcg+PD8YqGF9U0j8VAVCaWZJG0qlvOhWtKew8TzoV20UIKSJjPwyQt9R6BDsUx+gW2BZjv
aFNUzDCk54glGnBMVeUxcto9ATKvN+jRXBCPXV2o+3E6vVEzzI9NLD9P+ZLY9yGmCp/BEMWCgcpD
oxBKpoGIZeedu7hV5kcZXyJdIyEO+e8kUCsCjQJ0pKCTkoHpFSZzDE6BRZdf2WRo8prRrkibDS7X
qTpPLuLvfdN5jWY/BL0t3ilQDwESkHHDlGCl9ds5BYZyp8UVj5e9E4VxLBcQcdmdaimAoaHOatrC
e/5XA54HnhmQ4g0RfpmnuIubzKjjTfbu6/OaXloYahXwcMz6uVllH9xAWHMFCOUnRmPbBxdLOopm
2T7FhdT5E2A6sQSTO3m3O2lEuL7QFJYmMF66+mSbcaJ2E2JdARSo/GMqOhWjUD6/sBSO25NrIxrM
bkHnJCLJwAvwd5hD9I2YzwwsykZBs8GhflOQl4Ilu4KsTx6JQEVknI5f+RkghDGHr/UzjNCI1aZ9
sZO5vxJRULeXpLXyEQPoyX0QPJTDHIQ3Evq6Jxe3ESdRHYxztqPxjk5kaqb/+eDygnrDO3aTv8dx
9XNqCTbevmkahxI7ZwSkZ/grFfcvhWfqL+Z3mv/SDD4ydfVSrVcXTZnP8h7ayJraOcANFb3rvTSp
c8dyiODtoc8dIzLDOHQxe0sEZFvaNX8nhnTgLliEpgtvVT3juh1tOIuPUYJcmf6DVxbqZDvhvMZG
jODPHEcSBuUtxlGGIbfnOnHG9DyplxpuadtR6trGHmvofz8Of2sVsLfopD/5Mgj0AbZTAMbW1JcR
ketuwyXG4vEE+OG6Wj8d3Mb9ct95cXraJXGBlWhwGqgyPgUOlNb1CgqN2VCSAIDcXG6Evu1RuRIw
UWAQosc5j5ywziGStCjh7t3YudIYZxBgY4iGzxm47HfLNzeXGWJQgGT/k/GG03zdrfs4bk2kMUoW
IVV+8upyuXzSYSAg0ap8eB0nrcr5J80h8VvbC77ueQtinDVmkMZsYC6BEcujPjOjA3WMIn9TUPaz
w1Uur5ZRYvzwGamu37hiukoUN0I7EvLz0nFLMRnssqaKkWwy8hMGofoXTe8LY+KlzW83HU87gTtA
1s3MO1cUeoHBwnsmiTTFdJUjxAUYvKcpQZMOO3aUf8iRrstUznQ/u8Dbf59rtsYrFhh4ztlTtLjw
7dsKcxXWSNDzjvr3FzctIw7jxW8fqF9s3HxC7SLpPL4axXVx3nHt6xg/gaMxoLCdhgbsLKnVM6Sl
bdiouFfeAPADfACG3oKZEhKBDER8/w2Tueif3018I1jpmuUOjpIvUUnEdhsU1fQbwJnB+/ccxVYB
+9sexXWEcdO3R61n8ORMhP2fVx3ihp8rxtTQbDZpBUqvx1uivYbX2+z0zb9q3uGfc/APvo3/jXNG
ycbctidus+RefDqeOd/akUOj9AWqg8gDl1h/Exlc3gQTyZnFmNECu5UeXmoYM06C6Q/uOV0bwtYp
yMsnColmSV7OrmIAisoez+Zu1vJ9WZg5o5IhETMu7YTRUpu365CRpxG1GpAVmzlFZZAVGMNPfAU7
ct+giCjggFlgcrW1zU6IMwOQLpyPe1cupjDKRuFsT4ti1jjPJIJpf8zwbePnUcxJg9CCxZWxS3Nc
flnP9+KxsXxd+Hh4pE6oM82uwMxFZIIuIxQPzf+eC/zT/GHPLCYPLVp9oLEVebbjk/VqYKsQDGEW
ajz8R7GDSi11Y/b2J6myc4W+FOACbtn/jErfvbgNGHYyyeS1x+7NZ2npgsE1vl+fDfZInFguQ3/B
G0nB+OFX5cVf2JPJZNLovMLM1uyQVtShbOSHbN9ZROh8llHdtircwKM44NAqAIQhDeusBBz+jQyf
aCWECWQ4NDdqw39o2BO9bWyQPrPwWa1Fy8G2gWFOqVrXOL7g1DCijLsDgoGsi/FkrsDACyv1TM80
QV6f8w4Dxb5SRwtmV/3ak173bHA+uH8PCljDGgQYFuBwGFOqHgPoF2aUGJB4rh204wB3TGZIGGI/
kWFsVKOSwvUqKVwYGC42OlmjrXcowqP4Zd9zuzTFhAXlmiZt2bzBpnQqHX/kWxLACXPjMFuT6DrG
zfv3y5pCXhW3Kz1OPh6hUp0hlPTDe509z3VVAC8+q4V2Vzyu4KElf9R+HVKpgNrrgMA+U3qxX2TQ
tioamUhsajtmaFLTZVEjpetclIlw4wqCuQFNsfTbMKjVu+2PQIMj819dzLtSdrYQXREpcFeeick7
FXnNpKxke0et0F5YxpFzDWiboEnP6qXnmHX36fuCM933Sx7DwXTcP0u6jKhFf+BkGRILfLRUMNTJ
qlR1NCUQBJ+iTf2tUyczL41XP6R782Wb7s52KPTOLqyWBqDQcakhw4rVRh347WrCvVWxPiliAYMr
CyVTX/wV+owHZ7McZ2rG/1lMdEL5s1ngcbH8ZyUT/7KE5rKXk+E2Ila4439BfqCrsmEcLBvHbJ5Q
ppT4Pm6cYyBuYsrvQX40KY+7tDQ3ktq+xJQg24nJKnaaCgr9t8YXWv7886x+h8r1TP0+TEyv4Et5
OoMM7lgIeTlHAWmKgWoFA9/SkfzfUcXiM3KVCatOTRYBM9hPvD7oZUS8FedYdbHty9dGBKm8d3VL
FIYN0aH6/S+8XARzldPGQcyQ5stYaRWJ01b9+8PO8SMruVt+QmXWvGWxS3e5F67FrngShK+NktA1
oIrw47OlcSkDPwhQ8K+4NJ5Xty76H4w+1sroAzEHFD7rnkjfKqYbY2aY2zvewuj3w3W8bFf9r0wa
x5zq2iraYnLLeMFA5pqdhm6LAN+JGtha51JerH8weaqNHa28n6klSoZUMP+kEKzXwtAUEbLYYHq6
X3O5HJK3yqmIVjES5S6mebs99NX2fxtCQcudNgRYpe2UukuxPrci26DcSw6CHKd5y8tYB8QUtMmU
yZs0xULsnyhyb1Cl2pcpZBP00VmVb9Us1Yji2CQkeL1Sdb/eANIf8eDQ1E/Lm2oxjdd3Wd/nUh4W
omRCiKv48myclNIqI0JOufolxDle+bqmollho9aBXrVi7tLGSE37h7mro6XEM4sTkEafHZAPZDt6
0SCKroYB9JN6L5AAL4bqwfmSefpA4EZ5zbQ2s3vMHKXuSC8i1axJ6vxmk29/rXtJT8WjYIVMTVfX
fl/45ubVeun4muweD8WAhv9nZtAYF7MrQnqqby+uo5HqfYkFV4VTvBsKH0cZe09lWmuamQd2L0NA
P8z4H3cvGZ1HMsaIEKKWxcvYdlV5STeq2twDaqWX6mby219Q+vcj2Tmz5JDCxlV5Vp2Ock7iYEpK
ztRqLEQDD09g5CLZ7R09l8ZyU6zTSQTalx1YT+kaDcxSr1Lk0meykSRfgI9wKV9MhaBBgs94Ko0x
Xf8XcBFvCjQzZQJt2ftAqLDrQHpSqNujGFKYehL4Q2tgXefnvYm/RAeNpS6FfiCiR0/k2s46oRmA
M4H+egtx5bM7A7MVU9eL1Fyh6GKjQl4vbc/i1AMbzs9+UF2sLKpVWcODh9cUEci6MMPTXUub9v68
uqgCd7mUMcKW0xiktPWYLDiwHtnsO+xrR+Jrl2wPYETNaTI687I4tGzMwteZNnclHRurPQKMKLpw
wLG0Y41D8ZTMFDNcCs2MGGgrSRaQm9vC57UTvSYC+X2PXc7te7WRaUY6+Iky+ksGseO0lsDqWnRC
RnM4o+jREQosKTzm7bXnJYwKyCuC69xv6rjeTymkn4goivPFaaEDta+tYbpaeW9ARc5jdyH+aH3w
71g6oGyNjISzoHHBM/9X9UHDgUR8J6722pPCgwvpiFbStbPHX9mKOcqBCJOFLV6LS89Dk9kxXv5k
fJB13Lo6auaB9FtUkaGiswRqSz/NwFavs6i36XMrzD5KCp12SovHb/KW0H9DBoaTHnPfGhOJzL9m
x14KiMXH72UVjcPeMH8jtOA5gDW1RwJ3pAKIL0Vhll6IAYXwgM8t1NZTTkHNxPkqxTDWPkZQTOdB
XOl/oCLY9nlzuE2ICTvx0KeugTdY/LSMZl+v8Am+dX15i7p6tm15143cBH17k3Ejo5WRIdObjwCu
GO9SfBxFWvHefTZgttuoi6aufRPUVZsY4whu590lGfQ60Tq9+I+9ESqXvttwCF2ZnF0mJcu2VGro
K6kLjn8+vgprhTRnv6MqHHLkEJCeG0L1oD/AuPv1terP06vHZjlxNcEQL42PaGutphoCowBTP74z
fJFAtMZDnwK1h2uMTjmsMj7nyPLMj+bausQPdQCUDDiGvt8A8xtvbCH4UCafWryc+qoI1lYc3rMQ
7x10gJbojE/gXu0qlz+1L4j+Pu6EA4F2C7fkQuePVeo5h8MrJ0oHXtgqDogHNtMPKjiZ8obY/hOn
deXUTi2pV7Hgyfybnzsj8GfivcS8Ilsb+x/UmE9kjLO54LOQG9HqzhoEUr2JBm1L9vpWe29ZVPa8
LzY4/n0NusZZo3ETYLPV4VQNXE+RxWRvKxHOXPx0h40oDAsYWuGs+AoNISUJBmxH6Y4v+xBMI/xG
YZwKdLEDhFZmuc7plU0cXWFfs7/i6+7oOlGZSGlb4hwGDAZbSjnbTV7u4HJmk7Fj69/8porGayfB
g0AO6VNU2gTe42y2Xt4NSW+CdTEYlKPjCdveF7Bsz6CV5L/YGX2Dp1IcsLmBJ7dMrzJ66N6qLgoh
LvbhK+h5AZeDIKu7uqfio3leXuSTLdwGMQCDkwN2kK8aD4FO2JNjwEKUvH5q7S5ZLTWgKPk7Lj6K
vmb5vuHE0Z9sqNE0bxPld2DvXCx/oVaJoB6L+tZ6AmtM0OaCflitjkjCCJCS0VRfVbzomzsSYD6G
H7UA5MppF7truJM0MVeNeUBwsQxaOVGrI16E04z722Slfijr94eGnAjvCly2CCY6Blizm1AvN3BP
ilbJN4fEjAeexR6mNRjCBAE7EvcUbbC5dyX4tdUTFbjg0Ei2Fe1TmlMAeHUIBSOtmXUWH/ph6CWw
dfiqx6J666ePHfCiAnHVKzZjXip5MC06zUNUo0Hl7RcTj7ViaX1ZIKmL/F/9HW16pb+DjpbRWPKo
Lso2EmzhsQrE+7clISvqi015R3cO9m+3H/DbsIsPnqGhGzQA4+ShMyGED8yweUpBm6BurrJpWA/m
r+MhPjjFbY2V1iltFn6kFTRWJWWAsFhNg5Ju0p3maI8Veu7IDBII/uNvg5mBDUTHSwo2Ur6VCSC4
OukbacZkgdZpG6864rlRQcIiXRcppMfU6eTuo/6Q6XnCEtpyrMqOAvnmbXnCIStoFev2dzhMHRvA
Hs4X64aDGUREa1Ur9Rz2GQa0ZxyrJezUl4zU097p3rR6VGA6Gh2fcbUgLzMm9ekRi/hUfk/yN9Hm
+smP0/I8rJrwrOoS1OJvr0vRV49lyWCYkqisJmTvpWJGJK5/QNvbwcmZTwWdFpM24t+HcrCXtors
OCL9JeaXnrpA4797fNQ78e+wODlHT5EPKRfdHhcsx1kTj6bLd+LiJ+yDyLnvKtwSqJeZbc5krZE7
9V6K8kaVdsrmfv4K3ucqxHMlCzSGWEM67S/zTnwQQCXdRUy0+Fo7GkVDt2HVSjiZWai45Vo8Ny/b
iygT/5iBtiejNxn7NRwalXBXLaDwgMtVfeiTRdv3gKgJuZH/6NPGjKRCOmdBK5YeisRSh8T0d10k
CpJT5AYB2+DMJWAAnJbXjV0U2nG5qed92Z1leoILuW/QX+EziVL1VaAvV/i8hmpuZ1qRi31rrH0p
ywz3sSqGLJVAiaSJYb8ze1KijDSoDDeEYwZoB8Pmq9fDmlKdWAcI5mMrFHaa/Zn/8bMLSqG4xtWl
SDMnvtGpSbYB232kPFoTygTiODDGlziA7PA+wxMuvd9V8u26p1lj58X+RGAb1nw/fc/DQM8XDE1L
S7AdaDfeUYr1SCRoBlHFrTqSa5jDmZ8QvOTTOvEgrIsM0HB2k0xawrYftXb5ECTm+Fgx59LWf5ml
WWgeP/wwtRWThf6/wBW10UKcAOx1xegsHStPr38Sd4nPrlNuM2qacl6S/Q7LDhAmd9NFU61T+FUr
zqVWTHqqTKXYCHwDRnvqtzwze3gmfNjtBmS1rTdFNbzCeAji8uoT7ryiBuhaTvGowRs4Q/LYiL4L
rsBHuKaFdfeTJTSrNGM8wDWMxh0m7wbLs/+ZRhFgQ8/YfV87KAMxZXVEphCvSVv72c1Rr6g/VNRe
octYltk0toADv5eg2P6Y6tGn9CXdi2MXmTN3dQkXV/mppuj5kBFUWT/rSLSahCNDOzheIwdD92ld
B8im4ImXbqdvJsoz1yYGRLRt3wqH8P9tAlTKepwZgtM/SjMPtqIlWXcw5syRgKT35ESB10W6kHtM
MX8srn6nGgZRnm9Gjcsv+FVlPftBZW3NkozIuOCqsJjmYn7OFVRASO+jwTUNofTicwkRSoDRhfVc
CceOPgUR+FatlEbxvWVymtYQzSPRZ0n06VEM3zN6hQFV9wVp9BdESh64QP4WcXGojYNFaDBiJrb2
xnr768yObol/F8QJ04srjF/+9YPwfXrmM4iYtj0OaQbaTf89THyQxDFUUjYUAhkq69rUTWc8aV5O
XAvYxga0jEtb18x1j8S0EQqRA5tAue59Yp7nu1qy4ba9UQCduBeF8M9KY8+cp2ECy2w+NhueAanF
8XXoSGGZy5hJYgqYSKz2z6yGkvyArYQZwQd2wRj0H/mja4+CNgQ5ti0NqUbGzmaPSJjGmKh0AskS
QE8K9PElPk2AsOdkXejDPKQmUJk8dRWS4UucVEfnGTm7Foe522lgFF3Pv1q1BtFOcDjckdBeTkDu
e1K4yHG+1LrAiw3DSN/9ZUkgduOtvDCU7byreLh6lewS7i/viFh8HkpHFOxM28w6qP/6wX+m2lX9
T+sY8MWFzkw/LxpDC+pzmYtzYx67/01AnZ9DzVgAug4vl4K/v/JCCm2mvGLiFPWWay6nnA7Pju1S
uv5lWQqKKsnyMAa43RmJlfluOLbEt1q+GGUFFsflri5BjQDvVb7R3SB4b0h2TD66h/HCfy0LPX4o
gTrFXkcTs6kPnYd9Ig5IlB+VEYX42LBAhC0k11BRTrLLPOHXEtd+X+s7NU815BUqYCHBNAlWCWuq
Qpu+ZPh3Ez5e1b/gzfQ63564G1lIc8GA63ZrlV1c1nwSISD0dPr65t/24SvltNi3zURpDyhcJpJt
Wx4rfUqq6LbnTJAPvs0Ihs158ljEkB2shZrl+J1D4WXJ4dCMSH1ofqpkgcadK3aHT8PCeSmpWKDN
AXHzBaW+neS5j1Kp6sbb0v3y8I07W73Q3ZYZcB7t2dktAth+tzKRMEa1lYrHNTtl8b2noo1xp6pr
h+/mEfxH2QhqNvCrXXswS/akK2+WdgBCAGFvsgBcPtFQIMUpnYLCgGP3plthURWWrHjfABLbWIHp
fv7vwKWKlCpBCaUAb4z7OxVoJ4BX9xDeT6cvZK9CZ6JW0SmvIY3wPEB9DzxyZJmOPY5Qq1q0lqve
B7zAj46O8spvpHs9oiBAaOu+BzwIxkGm9AzjwBBlXXIssLGI+PNHhkW42+cV7HHA3wxqwzy35Gal
NvQr2YALd/L/vOCAhskHY7cP+9s1phGCzDPtVVO5YdQ9nc9MLuGflJym4dsXFneHaOJfttmezOB9
nwbiwZrVPd003ARVhIXFLS6gYynH84O9lemuhyejID1G8T4CXD/+e2J6sRSMgfrjZPX1rYyiyy8O
y9KE7O/BGruRsgQdnHmUOMKwnAnKtfG8lAhni1tp6+DB5rLcXEKnCkaKY4vdFeE8RknMfvTbbFW4
bKl36eWvTuUUNV805MbiaZIYYxSrdE74SxTWZUcPRBhBAL9tp3Az5T9bYPLoS+NL5SCJxVdEZNcz
gY4I8eMhtJYILaE+PoyIBejUBBe9M9dkvM65co4tc3aOjRvvf4BpF6C4AGgR/5M0fS/Aj5Y0g3q9
xaDq1mG/X+zQQFh8P0j74zu+Awpm9DlBTLfgUpXSxtuUzVPipIyr01G5ThVoJHWUPaAB4T07HH9Y
O7fMXJ2Dzd3owQZxnw4FGLyrBeUD1yB/Sk6YrIz2iEgG1ccPXhLyPU5YNUrpiovRNAP0spND0QyT
L9Gd8FeiGvs1seAebf1gHVPlzkZ1+fT7XACcEv+a2T75yw4BNf1hLXyp125H4DL+mKcnxmqick0w
wrWwfehrF1uyf49WvOyXtjQevvQHIWpCrSszh+Abkjf8MhYbjfuPb6wCPu42llYdHrKlacIvGOiq
ZrL0LgoBPBF8h/FgoCsw7DQinzx2CGu6HnGtHeUGOSYO3FYKeS7YjhP09WnAD3C+qAi2I0OpEdXK
jcGUgZoMWVfHX4LLcmnFNDyMWxO0HTg6b35om4zCfE+ik57dT9SK3S5DDla/eVrSv65Jz+JzVvHA
TwkM9mOqDicaxumZxy0BRF1F/JzCie1vgM5hLegZd7e3xMB0FTisZea5p5wsWln+iPbx6e2V9U3I
CzPA0lG0HZWwUJ6rwyTc3fDxh15ghRfD9Mie+rbkgDcM3m0uojqFU/3HMLlNZItVuYPubNLqaJON
o4OJmcbS6zF1BblaQLR8ER7Y2mmxB/4Zo3d6eKNrux6+l4iz0d9HzIfB0W0BpSOy8WTzTM/jLphm
4Bq5lwbOVSN/QyKdpqTlPVSDE4Uam1zThfTtOeFcu7k4Tw58TNoseSvJrpSLRCr2Su3u4BbdpTgz
kgzDVY52QTdlqSfkALIbBcKqIBtEb/gtkPbpdFASlocdNxBzsCqRuGW20SO+Ukp9uBO3cgSHRCln
a4y4pmJstxtaoMwQ/LWJU9JnzEfDBNNbZq6EraZP7YKbq0l7iN2lOnGIiaYHv8Sq3NcY2zyD4M9N
5oTpIrwdIZPROBdyaNozB/Rs33TDBUJOCs8Ph2fjI1nV6dI92YG+4k30KgC1kG7zrYdpqgb2ih6M
BYIDk75TVxsfCsA5ZNbtrqOOGiKdmPCT56lgy5ZAVo9tq6Ehw4jojfz4m80rllAH1p0bZ51CY3Do
0IfiIgaECQxLu5QJgl0MXL1Gm9Ww1OynYThxezaxp2EZS3y2dc0NrptIPra3ttLJh5s43njSZHDZ
bVbvQVvg/60/ftFVeBmM47adFKC/i4x+xnlGnu1sB9FE4nDgdMlkmd6gkWC2nOCkRwbcSgz9WHKH
YLg0s4AaxvBR10xGiIaFvOLt5xpHXaJ0L5mAZkQ4ELHxjeFUWnoAqNnBix7aL78sjthJiIBkTvrP
rhFI4u6t9WvXfhIBkme02HePYjXLQ/ZHBhT8YBUC9omDEHT5ykGIjGI7uC/dq//q1QYSwf2ljfPd
Mp+BeRnEv4S3oSBQLNYagnhP1cq0R5UpJfhTz0Cs9JrKSbYyk0PeFM9JtpI3+ysGcnMP2uheVO0D
Aw05xcsIurvsutfk3d3nYu8/XCT3Hx4Wf4HCiD8BkUXPGyenPcVwPfIbAXdcF4QNGlfMR3mGG2Qt
MLSwUHqwzyE8dCiCLIfSgw89kBIsHO9Qh4BAx3N2rJdaGnbGNMVVo9XMNC16u0v2rnFnY0c4Y0n3
fO4VZrUwO9X9yDuXlBUsaVsMSv+Aeja4w3OQDnK2Bo27nZWcNv+LmScIHl705dO5XIN+bXnN24Dr
e4kqZgOJYAtoIj9uQrqMWnv5uZIwIAN8SQ8s+GW+JWWC/7jUA/aqBDbDBCa2+A8LeEAJ4W+Ulfjs
gi7G2dwIT8+Rp0hUiDj8IMHXkk7rIEdxRQPhToR7X2BIfIUAflBoCGhB7Kpuvv5dk3vcSV2ZiR/J
OGNSHbfdpFj+AkS3YN+WzdMXlgoi51Y0okQq8urOLxDdl5mvvKiFw9DUZ5Gjvblk5cpK0p9KvPYf
PCdfJyJT1j68EgDYF1GI+ImDpoKvDh64PvPFUP9MhMpH10iaTXqBX7Cr0IBvslsENd7tGNThRePx
0Dij+6i6+U1R2jiDYM1pJPXCS+JmBgS+ihJLqRxDdpfPD6NbUMfsmku0hdlYKj1PdfLs3SSW/obd
SLNAsYyGkgkEL5OoaPVTIAuGhOHPag+11e5/pSZcq849oIufRDq9HomIAvZUiyBeos7H5kSi+f1J
q3qnuCfD5bJVG4DumhYII67+4mrgFSBvLr/Q99++wkNdXNavv+fa3T9xIKHeif9Kb/LIZu2h/3os
+xkJni+sSsVUYyAD9lMXVggvnL0esZIWpEmuegv4beUxMzoyeucvBDfnVZ7mKdmxuVRXc4UVSwcl
/m8NdURl5GtxAeNqkZZywxpoliM4QQ7ZD8dBo+bU1TvU6gJ+Rp5H9x/v1/I2H2/dHK6qZrZ1JZ3M
qnBfWV6hUqrqbPgqm/yCHCh/ABdXgOcovIHVDhMCwYSXBEQlaRPZVQvraTnmieAM6hwn6PKlGrxa
62zYtYdrrfIcXRyebYoqdSpkaUP0gXInWIUaM4cFsMOjlT650NOR7l3bAxBUy7oHPSeGxleUY1BD
XSi7AYjtE/Xag2hW9NxP6FGbJCFJcu/yVP7y0yMHImW45E7YjnfmJGLKTpzD54XTWK4LDSAEQtYw
7qlkhMSlkznvP4vgrqcnxRU+Td7T+DFHL+3guzKPnN1blOHT27XDQ0meIt36PmkWCyUV8ia7+p5T
y3DHn5TX92nMC2GcxcjtNQlWr7YS3HQsbPS/NzrkFoYhAnfsHWFoO0LnfWQuwlWN0ByNiVgkQHzL
7VsR1Hl+3iKS+yEBB2ULwrwSOmP/HYzRR3DQ/dE8DnJ77+WJU55VvDRmqwbCdpx6EEBn2GpEFrFt
6XDwoudrv1w+2R9ah6WPQRunZ5AFfNC6vBtUXjFD38Gh6dWYgb0Vmz7aVnwcvYBcIaEii2Vt8Twh
vOYs/ndfDqe37Z+xuu2R+7W/rkLPC0UHFkD4iFXQKBbSu1YEA/o8WK69LV3JaGfsxlwbvm2rGTpo
ioBOJcTUoFEzHH2hefk6F95skXmsL/Dki64pDUCeejrqvMqq+Kqbg8hY1XSeTIfq4tuhObZELzL+
Q0B39bw+PlPT/Lb7886Vtu9qmCv7nvOewQ6q7bSJO73NMP5SYHMrW5FgqevLDIQoiV/SbulSUJfn
fIod1zjlY+d6YmuUeCi6JVB8IlOQ6K6K9gdh9wNm5gD8bPc9LoCEGfNQDp8R2XhPCieAt2s5Sniv
iOA+z4X7tAW+g3oAFybvf1v3NwjyPtZXFaybViythBha3sxHMZLG4m7lt3JXCwgKlxUO5UQCHcjL
JPVmS5kwxnOujJNaCBcf4vpJxcwwZzBIJrx53/YKJuGgA9FurtmXReQWL1pmLN+D3nG+xmLAl32p
JOgL09O13WMOCtrJV/5gY0nPNrf5CatsPKkGuNuFG+phMtcbaqWmMi8AIt6juoV8oaMCR3YdMaNz
xtw8FVoIXQRIIngcYTrmjqcW6s2DvX672N29NP2R+Gfex/xdKo1+gRDU+DI+SK+jw80EtN01jBEe
zVE/Vr+YqJ5pQ6/RDe9DAKYPFTJEJfOjlrnMlPeM2LGHjlp7SjSdjqwPpA7IuB1zo3ehctVh8vDo
/MWIIxSp+NexvQv0r2ZkAb7/BQRH5iN815djJF4nXZv7i+WJj4+B0c6+9hdklYWUOey9Bvi6atDz
S1wpUwxSEmr93LWnEOL/XGSPxxI98xS0kHo3h5Pl2ycGkPILJ+xUXLvx5QeQhJkMgkSQ0WmJTDTF
GLtEzhYWQTeAsJ/wD3wcD4U4l7c9oZb21eogodTJNJQDAbZGf05YtKq8F+OhZ111uJDRD/+wYU9G
8QwRTbP000OQooYRQwCLTlDwDTV9xt3q3Muo4LmcWOpYXS79tgRrvaep+ocjvCnt4hMROK+tElIp
Jp464Va6l8F0SplZhkuhl3IyygV5k/eN+Kx3kexJGFt+qOC2h0y/RHOfDbfOcnI6lO8HveOKLvvJ
VWlVClH8ahtyIs+17oZhQRSRaRFesmq1rrjmvL/8mvgbHlfAbN+2ird4D8LWO+JYkae7XY+Kde9F
8ioZYjq+1oHpIrwPomRH1qruIfmsNOdSvJub3sbD6G52zoZgQaIyxn7pGz/zfLP4epVucwFxxPQT
pwuochd+JDXSq178g76chnB63TyYwUKV+GG+9wQdHjmiyHrBGNKmxcUGJJcjAL2f+jJu0rU9neeo
Ug6VQgN9AHzeZbA4ybKgIueOHj6LbEGhFKzPR2x0F3FJH3gVOfgdoRjLQFzVXyRAN1xh+a8gWZAL
QO3TrJr3C1j2KTu+RSW/5jry23Zon56toKew4vActM5D65fMOLFPAwD/EWOtV5q6sSOpWWXlwXNK
Q5cOPKoqav/dzVwumZB89lCyFXLDGzYoCpjlrMsQw9kn8s8NV/yJHWYkJSNMlmXNWepXdlhCO4kP
sCZOydmkP/OQbXkDJzx1muxBTKBrQyN7H284qDu5JmjKsork3SHjWmrR64WmupycN36L0IfgSDE7
41rGjds7rOJhLgog9LRfu9SfrpCxu91pI2ApfB5yUK7VuEJ0Gweg648lHieSUVG19Oa4Tz94iN5J
dRBMidISWP+0jjVAc8bpT+4nxBgRxdriwSkDuN1E1OBIPFyslBy7zBccSpP5eol8aDuktP3+jLsN
B6ZCp3xJtcj6ePtGri7iGiJsYiW8MmGdI3TQS7BLjpPfx+27UAvJXs1vqPGmGpahM05CFJUnpKG5
HD9GK+PDPaRULyV0vPW35H/G9f2/JcZrZkrnLFFROpcRxnHpWN30zguOGOX/430USU71RnUp9hZt
Kxb5iMyULhUS/8gQvQYaSycySoatvOfLduXjQOk4akn3V16xd4eYQG6/UbXSMxEcCBM+9TBmKPnV
T7ytodEXifPmX06dnoTB5pnE4alORpAWLmCn4AsUs/Vs+GBcflWuN4zkpGE+vl0UhZjCTGbgwDjX
3vyirkiWrT1kaA9HtRZu7mUX0c1X5jxLsgCtVUa250ln0dUOFdjPPBWRvwbX91U6Thz/4fz6JOQl
es3lz6gQFXbyf7puklVo7bBpmfOQBaYqVAvc/JxbUO9P74kgQzXxy6DZcPc7QUtZXijyIzGA2pqA
MyV1+82rb65NDF9srz3TtYoIGGeHFT6ZZSQs9EGXj8xIMG63SC0PHGkFS3gNCEkHFxVFNGhzaont
rMVE14ZVPtGQjCkdcg1f1LGsEBckDQbv8mQPuo8TlrQdyILvxbQ1O0QYY3H+9WekhSZPOSaX9R3T
hEV7iEOlNKiULFC0rPaaECMKpCZauvBhybmnvsbP8Dp2Zn2cMT6tVHowMkMGBGztEEHBWcuCFUen
OKoT5vxWAAYeaTYHuoWjtOajgDuzMCqeb0HL2QY7d/yVsrei33FdSQeyYJBJPYtzNfDPPsdz5bi4
gDJb2XkrvH5D6g5vRGRiigaQyxG4D1f8h26yk9efA0Yto7tsnqEiaKsxQdM+/fRJi07a6AEl67YP
78iviD3qT/PF6vYV3v6xo9QHxFa7Hkd/WfVoQzvfZZOlIui0VrqXedrkYruihrMwOkaRw5Rnkqyi
FHVJG1zarCq7v1c/EwRI2kzrj2/ia3kiEtu3fVK42Ed9mbnO9eBlRgGcBISc/3dXPQkeO4deakMd
sBFBIdOv/LdT42oaieD39KvMQQRr9woQLeJWlrufrF/HhP+mnewkDftz3Exzsk40uuuZulWe7bXy
FG1JIbFAsKS7i/u8XRcMFxk3eXP1a4F3ZRW2dTqv5/X/JS4CpkMR7Gf6oDc/ei251ma8/V+FmIKv
lIVCei4/HXQNKQOI4BP/+FGr7ORDtpYUBdN0u98WW9Po4CJK+5hDAaM2a6OISmHsUABpKmAf9LYD
j5YKuSHol/l4ETOiLHaHVY/uKlqUydA/p4X7eT/jQ/JtyBbUcGtlNaZlXgKSp+C/lv1dtRmV/ooj
Dax5gU7kv7vau0QNvrcFeeqIolBLyLqtd52PMr91GTmMHEdgddVArp3jJ6Itsynk0iVWUHN56oB5
Rt4NJtvI8oBtZ5wMbtYL0yExghBmg3ASwH3qXczcTRxJAYBjfse3IwbF5xiATSsoZ8B72SqYf7oz
R8/g70wRr72zsFZQNAS36liHPZ9V6nE4RSGq0lrPETPmlrzXLYypwCgdZFk6HxSzVHCA9Cb5iH21
Rb7ezrn0aDPNalToDGX2RONEv+U80WWB03npPhRaySeq3PcubZ8nxzyqgtYjX43aeBccycaJR8n2
ZbRmVZfNvdrffkL5ua1eh/abK6uHH/X6khZuDiJmTzG/AjEA0GINJgxNN0F9urg4dOpaSNRhPqv8
NPX5uzJ6/bK3CmFRlfIZY1el4f6BTRSaak6Oo168d0zQ2MHXgGn6yIt3vRuJErMdAQMRBFuEXsZx
wiggAyoiIyo3G/ijCpXLpZVBvE8flRaPFZIw3P5dJSb5ynt1NRRuIk7zH4P+E7C8/BO7rOoGmw23
FaR9A2LpMwJBv1I2U4JIitKUIx0VSEwHSvxzw+fd/OtgMok/ujqYt6d4l2szOE+Am9aFxvB1D8st
LmCmrSSN9C9owQe8QcO7tTpaPo9hKD0YLBS2kUHY3KtZ2+/+SS/E9g99+oeJeeZIJn6p4H/ZLJgD
h/uy8QVquzTHiyHkomWvYo6p7LFw82oQkBskADUQhMgObL5Fh4X+WGnWJ2GNrxZJ92xNzu8qVtG0
oLDQlqBdPnkNP9B490SoSGqW0wzLPkeumtAurautGWbd9V8u2lS8fzA8jgx/O+JSLalltY4NOSkD
W27YD5yN1zkdhCuEsgMycKC7NxtJmv7osT+4niGFNk6Xwm37GXe61CRHEhi0lX1N0Zi6VbdP1szm
Q3Wn/Yg92UidSVIQWzgdN/akAVZQn27y7DIWtWr3pxmtrvNssNuMFlIhEcbdvesh3Uj+X5pQXTmJ
jEs0E/jf08QP4+UzKCjxdggdtGp3OPhfzhSk++cTDE/FT879fBBdzJmz40riXX2wtEHPguYHUbHl
4C5SFH/Cydxqbi27wfH6s4i7eTFOzvDnrYf4cj5mbfGZ7nBFrr2MmIk+GpKiPeh0r6ZJT2SDfpbv
lYkkUYyVsKfMkJtrOdwDyfKjrmtLjv1Lj0fs/5/pXo2uedvixq0I3FsyYLDiMjbzeKu/zg17bavE
gEGyu6HC2POT13+2/BnSQYe3N1eQmZKdq5Zkb3zoqf2OEGYGXQY4IN5rdb+OERMEs1F4+H4HPSg+
mzHRwXj8/PLvt1sWtFtcBwF9rwyE++23b3bsepXAeSWZhL0/DZJCl5ryJHvQSVewFKRW9xKkDQxe
OP85iNAR/k4kOTch514yMxxuX1xZ8vpE21S23FzMYxKT3p4h/o/Wc/nWcepsR3qBNscEuIqtOy6L
8iCQIR6ddq3Fy3b3O3e5J7MpQiCsl9YwjqvqjPEyM2cIQ0/gnkFi3pb1InFa4QmGcBxBKPHz541N
b2xH+LEBz1id7UYVcVq0KYoVTzWvg3G9Tqxn70ifkmVSt00VoLL/8EEh1G9Bj8Wowb3Khxb9DwRo
T6Z5Nh10XfPUsRxcPKuAik+n5D3/AiNZV4yMphSA94H41F8lAC2oFFmk7IWnWp7kLsb6/9Nx9M6V
FpfVo+gl1JTO/9dII+Uy7d9SalrsP0wRPBhDyQu+UFzsgABNMpyRRp2ovdkhiwOjMcCO9SfA1YBM
Ixs6m13UtXzPnqGtIr5Kv/4VJu8yF0+N7Is1muCPHacgxYdineGxadcEWUNsrozYa+NRRaQx8AXK
Ucn0JlDb7m2VB8fiXuQwlgXAEMM30t1EhENBf8/zImhyn2VHQ5ErL5Nks2GZS7z2JJnM+643AITR
jJ5cyrw9Ahxy8r1e3N7I6P00PfnisCfif8G8kZAhng0Zy9zhnMImZtxi1SWC+i36msuRQ3Bxgqwy
hDBjLJpH+UHXrzURCZ5tzVepPfPp80jJzywmVUlWeONbUNjkmRiOUfpobt/EaIj1TforGGy2it5A
yxpHwUgjIsN8iRoK5tcfHJB2Q27SRC3ZKZQ+M2pS/CA2WAOf8umSjudEgeBBc4vfF3e2Ml7gIKyz
Bwzd8qnTTCp95Zo1HW6EMtWxKThekF4gzwxELvtsAFNbXS2TAnpUe43a5k83iYlbGHELUsg2ib3/
eMXiJUCjkJkon8uhf9ZZDUgpTvBN29ILHUrQPC3iTsKTgyL83FePius2xdmDu7bloMYaxWElCULA
IQIv8G7/SuU0GD/BUNVYOUdZEiUBVO8qZuP8MNkR6gflsQ3rgVhaNX8C08ioCq5BHpYPlR3m/W6v
sjHIBey9wJWKwPyJnGRRJ2d2cZ6J+RpLPOXS2titSfR8xALpJTLD7A3yfZaN/wRp1Q1ggOdwLQHn
jkfAaT7djYQGIJbYY6A8qapj1Jbyc+OhrKMvgEW4FxIWvxYxBXOo1QVWFUDu2ZwyXX9TKzBGfGnC
orzLbBfpDNi8Ksmv6u3h3cC1MFrHN0NrdEl0m2IflHxp17XKSPFAKAO+jV3JFYoDEobUIafTf3tC
EjzL+d6TIOort2zmeTridSSE8vPo0+HauUchT9IZltFTlRunq/cIjZ0WduKNbOsHwSA+2ynWfS1H
RliZq/sXrgkJNtP+Io/RQE1ri+xU/VjURQM/3509HB4gvjRbBkW9vNnC5mJZoZOCRCyLyJnUsQwx
6mZGf7gJQ9H55uG23aWi9nSHPdRWnYgl+WYo9JaYq4g+X7rWtT9/46Vcs8JaHcn90HQj5ggwbj15
pzXnWp4YxNYjxV2hptjmAkIttJ1peirx0KBG1Kj8F/x1dRO0qyfHZH/PqZIvnmlZWr+0zN/duxt3
OmMP+Pd8DiyzaiVi/l0ctGkKdVUc8bH6htz77/qi3Wy5bdeu8tR61B50me3W9PkCtsKIQ1pjTmS0
G6KsSBDfhOuUjMG9cub6WPo1NlqDmZynCp6TQvvyvu9R8hgnNNmNXFjTkEFIRLqybwM8mzrlsRDs
oiLqKyRYYN+JDShmwOPL39dh27aoQ+nFZ+YzjCf7booW2eulbhekA/3HOr0orqMIDGK8Lrv+J32E
PiNf3kUKli7CG141NwhX8xvZ2/v237/rsa4qz39+oE/GCesSrPSs+0d7XVxNxgwALY6OnNQx2dz9
atwjzv2/u3obzs+vcR3zuhqBMwYtIR461T8WQeDkAcuw49oBGyZJb6BpZUQQJN6h4NvAn7eIjVwX
rQ9uAUtMFxQX0VD/LRcGsIKI0zCwxj55B2nH0WT51ccggR9GdNWKbfSlq+wZu6iYlQrWjYR341QB
0DxJGfZXBaVxuj69pmj8Fc0iTT+94Ll+IQQ8N2YhGE6vAd0NNZu37AvyZ5254HgZUDERBHtmJfHC
/VRKI8IL+/B87+63G/2Vnwrt1wcqD+jfqDzth6r9gYN3WpNmoAD4VhraJkbU+dEvAkJye6/qnvkP
aL6KHiAhQucTdyunxM8mUnKEzri0HdwvQOoIq1w+6ydP4F9l4ZZ7zwGnjpXAobDooKR0BqtJWgzZ
vBJd8ZwVpNve66OunDrsCLRy3NfK41HzcE0EyZ6SCgc8UBa3nval6IWliSjFAjRKGRHAiN6FV+qV
/a0OvbWnKfmJhJXbr84FF2mqEbk21vhJXtWs7fEdRAWa/XbSgMX3Sl+eziNHGBHwXnLDA4VwoQYJ
PDQgo/f1CvJyTqhtkqvSrkhBpUImvhWR80e9ReUUOnTRwyQZ4RC5/jhnFWSiDZ91080F9UdztODj
CuVtaEeGpSCmv8vLu+lWpgNOs7O7AxCDbaxoPgy+9CHEQ7LeZb3qyhdizq6pCmZ9iTutctXvysVk
304svXu7/8Utp2ChgcygyVeGxeRg1wipAzYXUiZk+VNKNs/U/A7dbJS6cR2+pJM+bcRxyUD2yNge
8HMfLij/NghJMfkAm6rY9UFgsMWDGmwb0gSZyI/V1wworCENVLSsJtlbXOfkzpO9qoZL936etXxc
+3wgKnNnrut7EFgSW5hWGf9iXK7Tq3AocdDuuOqEh1Xmg/Mth32u3GN0/mEbTXJTFaukls+T3QOH
qyTGHjIuzSotmjDw3GjIYNTr3e+FrJQn56IGgTXVulYrKaVPJjDNltzXlIIjP9GFKPKEhlVGOdtU
R9gzpKU68vyPqvcqFU3ak7175NdWaEtih7KE7Q6HkYVpeG2elfiO9QUdqSw3sqTjrt/drvPehrB4
ei7D5XHnk7dkzKq/lUPxyXBZ7roopMncYk0rHyWnmLNmMY/UdTlw7x6vJEe1V4YaGhEfmzQFIrPC
wPJLkWRI3TCd5ReY7yMLBI1AWbIEKyN0jXMW0Lx+jyoedEwdr7Gv0MF19dxGOVcv/tT5F2+kpHW9
bE1K9sQdV8u+ADhO+QEQB+RV32Efy6BTCI2VOR7bZr79+M9NCJsIxymR92dQTGLH9RYI2uufpsy+
f09dNQfatBEriTmygo8ZjHmMVZTUgTrkNl8gzBfAS4K/d8tEYV++8jgB3HGjgtdk0UmUaR3vjyFN
fvdWdFCkharc4g6NLDSr30LxYidQ5/x+DhhGuvPdkTXA7AJmk9S5d6sS3qK4gztaD0q7hbdUxO8I
J1576WHVfZPkU+ZXfrCWG/f0rACxTBn/Jq/w1LWaPtg5mryPCcyo5EhraJXmgoxMXVKD8uZjyLzW
beWMN4+YLqpRPx1Vkaq2y4RVJP4kbZHTwhMdlZ7NbjSqjzn0v3yBqpQthoB1dWlBLHmfSaTNaV/1
2+9Y45RG8pYE9V/7gh8R2wsXsuENSeBJu8t8RXS2BImgjFie1fCmZy+yaBa5GZpPLbxyZhMtZx8c
A0w6Iz6rSFSpO5NvY3AC3TvlVNcxWfSqdYRWSfWGFfu3TfuW3KtSAqmYb7PWKHiFdNfSimqaCp2+
OXh0tvT1VsEChAkzhnD2uSyoDtb/QbHXAWo5BGnwD1q35e3gWSjneiXfWZB4I8653yoAPpTFOUCL
5CkDzxBreKkJ4Zsvtm6cc6+iuTn5F3325AJ/jjGXSnUHgQgnW2A3V07COc8MocGWJkEOyBC+XVsb
Yd/Rzj519aO20jPuG45KFn5f1ba7QncTzYOLlA1WjzFA8qVFVw7uRBexJ54QOPX6xSSGKc4S9SrE
fHaXEanZOBnWi/BRO8YssutJM7jiddYax1YwXBxL6YBXqtmA4njswmAYKLRm9j2usvxTytFdqriC
RB2LEPUY11K3ZeeNqU3mYEfWjPjY0DVdISDOTAjng4mO9FqKTuQh9PiAb4hxNojafk3aAXsIMS/W
zUP62Ysn8lTgWTJDXY8ISUjCDIyFGTScC2M8kdj1NVpEcoVjgHO/CZcwad4hLMwAJQ9WoaEqXngH
SHcHlQs/HZxVonur15GnGik4AQqBdjHVBI6uJr2UlSUP93lJhxmyU0/LT41jOUUvbKyZHk49XHhz
hwexPGBdyPglfs0ysZ/+Vcfwcl0uExJcqcrhKXhgCrKTtaGu23Ed1n53l3F3+qtL1Fo5iUUcYfp0
zu7XYjJ+X4VDDV1W7WsPckq7mq2US7H6tA2QwFLVyKO1jS4q9pv/KOcJYMEP8NEkD/p+4067IwrN
yT3rrAawIo6lyUA2DX0YGuEJGWvABzIjT/7JmS/l1VMqU96sKXbaXYARErLR4K3UzPyXZ9vy3Q4f
zvJILCzNQ0HeesHHn54Yt/GG+Ws4u7rGPjFVTZzXkY6IuyQ7XNX6WAeSuIfEYI0fc75E/1+WlL29
friIFvGndkQ/xAq86Fn0jXtIaVDzrzw1HxVVik1DbasYNz0tmpmbqGVpeaLT4qDVIfOr3SR/z5Xm
8aaGSRv/NlPx7BaQEdcRI5t2WjbkSh0DMtcokorgz0KMrIyTx9KmR7KV9M6HYbR/mwNzIJX4byC9
TGJTiCMu0TNjVI8NYju2lslYlt/eBC5r1lZN2kr/8FApvLZAlfWy+Ly44qL6Alp20OKT5vopE/QP
MgMOJUcIqkc/dRouGtWfAb08y2N04nJgyRbDFm0D2F7zfFRsfUJI7QI2EG04CByiRg5jhkQ3Q5lI
+x14QNPRJMjHb1Glt6MifBl89yCttxSeEcSLFzXaaJo2RiU4BtmSWCoIzZ4/DLslHxWtzaFV/MJc
SQd3ZlTdXlv/FZrwmBC/P6ldxs7ro5oOS+VJgRK0dyRUXEY+iGVvZ3uikEnDgmn6iULBmmwEzJdd
K401TX/Ch+NjOeqXeyqpA9eyFsAJp5ewWCzTpxj5CIbU1UKLTQgcjSk8aAAk1ivBIT1KJywfUDUO
ANSkEKVfWESJIHtq1z5vrqtrfcObeh9KTKt18KoA8DOLVe37D9TF4LPAOYj+fgNmlCt8xq5G0692
ses0VEbgMxnerJ9BuaVxHnKXofgvS39NZ/F1EZRsA3taRh5hiq6e+n13Zm0Yc67NvSTNlh7PnklF
xahW/rHYtazcKrj60eSGza85gpudwPIcNiLY5HqJWRGK13ruQ2AKahdqddGjz9Uzyg6HJ2ssuaI8
O9+Py80ilQo/Nsw54Yi37jLnI3HrRphTpL0/Qn8y7byTJTzONlAvFCf1xTrPyHQUe1QBk4aBitsG
cdCcIvaac5dOCm0kXK5qR2kbz2jcyxL3QalZHE92th4IuOXD0siIfCvYZ0Nnyto1u2yZ9bYXZA0/
6dI/xta57OPYp4jjUYGi2l0YLDGQqb5d2C6q0ojIYbQfukFYXf5KXD33IMuNnYyhNICMAOfaBScm
XfVchAtB6oHQuysPqlrOCCHoztQiylFGc9fVFXnqM9wR7qnYO5WGDYY1OEf53Sqx98UG438HdZy/
4jbfrLYy6vuE/8+5YGOR04Vtzhk9p+KxBTvOnSi+FMV5aDUd2cIk2labYV5N40EDB6sVAPBokKpN
M3o33OjookHNySg9qs2jXuaNa6WHZoRuCXh4GIH5vowBIHAE2tlD2PxgUvpS5/TBhywPmug+5j+3
X+mM7gMxtSXGNIKxmWhqAUf7XciF0g2fM8N40UuOUCzOMDRFplF8BhPs1zzuz9q5YwONcHCU6yXi
sVQYQt/ofEVl994bAaHe6Ou6m6kaNr0F05jQCNNDqNgxhXR1YRgr0hHqLArIZN7/17Vb624/SsW1
8fMTsusDvMPHWMqfGCRYkoHCr6+McXREaqg/lt9ySQzUVD7cuK0dbsVhk6h2dvGVOwL88E5UZ5GG
zmlyTi4UjT7cxaJiS9FUFNhFU30OZtDwiYsaKvSDMMm/58zXPVGusfApEP1nQQCil4wsL7wJbNd+
xOOilQA+iBjfmBMFECCN0r8zQrBtDeUOD/x0JolHFHcpQxHAqkBzdbCXCtQQhGU9Z8m4APf5LRub
5A2xNmOWkULisSjXqvn9zg2RvACBhd4lWPUZUEg0v81Ghos++SlqshSgHh2j6SXSR6N38jXmlRBb
RZ3SvOQbO+HhH+5J0OapDOSuJVuP8etnc61XyUQo+Gx4gIG0EJ6k6CP8N+jnn+tLK6KJ2bF5KYCn
7we7uO5IRu0WSkA4Q1nUJiUSnuUnRpqeN9Pmqg3UrkssxnqaCvpbWcNn0OY5Fe5wNbzF9C8WWakH
dOR/ZQwOM9z2so6+jS7wlBV+P8ltcIiEFXNJ44P6bH7rXJSwPvR9spZT5DwWC2r91U7QebTzR+cT
Xm5Lnf9SR0114aMQYcJBveCLZSTxEduhmtuXSf3HDZ+IP1Q9oWGeQFeW63lSxvpU/jsM02WwkqrB
rq5M3BEvV/kJBLQqlUsCif+4NO2Il6Juc1wjEbuK1130L8VND5VdglTz2lbX89776kZyaqufAmFE
ZbpvCrTOdeC6pIMDbRwuDcXQqOEGqpezw8dm1LKSAKbZKORFtmSOQnGsBJiPWWn3FH4bdxzfhfPX
WR9vPWy9CFNFJn57DrIFHxRQs4I/UcVmwNwxOrwm6S7q6BtfuJiSG9rgKzctwzIrWh/f5zlDGgaZ
/WIyhKkkuM5EqnC4DIfHkSy8YGvsrexFIUMoLYNAy60yfWtWFYFLqgJK1GOLvPDXFus9L+m7/4/m
5v0Nsk4khW6/pdPaZEwSEzeLupW4AtQLjoGgiJjvAlM2+K1aMzICRog6MjkjQUCW6xzoG9U8Bidh
m3i4fDNkQDkIKXLbx5zboMPnutpLfhhhUGIGTwoOvaSRTCfwgNEBHfVGct5Qxrrg/vPzWnKUPN8Z
SZWC4rBjRY7yc1aqyDkTeYGmu613wmtq1bnrSWYEMdDIfX/enbWhiZZxDae9Z+h+nzwMU2t+45Wv
MCswXHscOspkfoUzSgpABSKVZgCdFW0DV2l0jFZHBe1ab6h2/daR12RxB6tkLwZ4MT0DnY2AJX89
BXaLRB3JvZT9TgQnPsuHlXf/10ld2xa3PogFOFtyeaq50lRJmuT7YJxHqg5QrdpVn3VRUVfHswbM
EetrCxh7pB9Boia9p4s8VhgNO0pIK+yh1bB05UPAHUxMa0l/JiB0S74Gi124mmBHkBlEWmQ6SFxV
azWWM3evGnwrinNV9xxesqugc1c0eyfh78lyjfsCMBrxQT6h4pX+dRFWm3TUM+WPlnB5qZmFgjCI
sEr393+lBIP6I5nWCb0c5qE/rRrcZubTVyTB5xQJi7VvENgjh/mPd9R5/Alyn4KE5d23INwOy3fW
QH7rOTUq3AbeNsEwE/YVgQ7M2cFT53fm06GkSy+5M8JGptI2U0ADb1dJ1YAif196VAtRftZhZZdj
30mDgJ5yukSndfis/5uhSEUnCJRF+XnGAjtPtswNSokRJc4ka8G36hvcYIC/WdnrfZDyE8B5DNzI
tbrA7g7s4Lz58ZS8Cpx7PRWgJxHy4I/q/K68fdvBIaOXw5EZLWmQpgSyClLozPmuOCKGLcoORIZ0
Y0TJcg1eNEw7njcuMeibJWF0GxmIypqhonolcEXA99BPw5zL5pgznF3zrsDdq3LDRp1YwiiJuuzU
70P0G1HIrRi1+/La6w6eJeGMVAo0XxgIY8sx8NuA6gADT/t5LG5cbe+CQKrVVEj5gNYwMz0EPYOq
t9aeQrZ1Ecv1d1nChWRdhB95xHgpbeLDCiEXHz8OFwX49HK18t+8aFi5cHzTxFiqHFqgQaJ8YJlC
Lp4c3MaNEWRMUU0L9Mf9F3k6jVMGNLQhmHFHOO34Tw87yWNwZZe5cKKDeuhnxAANhcM+NE5zJRYt
a99UDGfACH9eG2UW2fDCHrWzOhc9xbkrG50kbDGKJs+a3GFobid/ZdgrptJ2zcdl6khu5mgqawKB
Y/7a9E4DY3IiDwOviLZizhLI6W76mG7h65lJv77eRaX9CfI9flYaVwZIOvg8MA1ijBmYCLZZv9fY
cO+wnzLdI4JlvVM6bLwJnLj4d+1M8vmvj8vsRgDQSmnwPpNFf8fXu2nh9ctlOnaI+O7yOTbtP3ok
fmZyDbHp8Ak4hcgkMnQYpR9HvrWF5Uw5lPirKGRp3fRrGQBwFUhw3wLD0K+VAm5lcp0GRGdpTk6J
inKDrvE+ysZBtTdLh60TLD+pEay6suMlZI/ggXao1frcWTUppSPYYHgdgrZArjABiO8+YKbLhaki
Wrow6dtmdZQ0oWOS0QIgGHZsPC6AA7GFYy+tSqsHHS4wGYmsPp6fYMQwPXXhVyb4ZGGxOVuJP0H4
aZhTfHgRCX39Fm66zsno1lIycjqw+U8eXactpQv6/MH3UA1DEE9mN06EpgAafO0ZxB0zQK52zCQ0
I02ICENjFAQSfWS7dxmdHGK/PiCfOzRaUtAUgsdbhm/cGqjdCsAV/k9mxQsXS2V1L77o5z9sdCLE
JT3uIhF2CDwrwxV04qLAeHYGhFXe2ui9mMCej4G93m1HZgEAQDepnLYuiexVFvdIgGsJw9jPUHzL
SOd4o2YidWIvNPTUOqHXSbdMIBivX/EetPP1nYwpO0RSot7S52hG9Fh4XEzb5FiVZqXzth/Qfl8R
M+F9E6DkUvarsPD3ujzdYERsSqO2C/TrTvgt/SFySC/9aL5wbbBdiPNz76vKYOOvL3S3cDub4tQr
3r9ikmDnjObM3VK6LIuEMkWd7eqF0hDTW6LS817vjn6+QcweHOz4wuhW7FiqgTwXxAbpRDt9CR1b
v/e8QmlQ4uRyEXBSKSvfzQ141oqljEmbFxwGje1bfQQk4u/d8JhUt0xhg8cnafoMAcEXru60K253
MuP7askrDjg4hnyVUVa5ECbOM02AJQ3C6vFclra6O60r+Cg3/BfkNBTqXzkEe/9mS+tXSFTmLU/w
/hoGnyq0Dpjtx/g4IFroRDvhxENPKykYt4bygQ3sj/vUsyKdNWAQ4U/Ho9QqTPuTX9XKtAUeGxrL
GdiWkfukDNjyzIObBYb4/pRPmDCfJAh+SDh3nqUwFuRUs1jBKnD96UXvdcw7tmeBnjeDKpHuVIym
Ix9Z4xA4arjmkFG8An8JPwn3xfXC0sNhLU03+tQ6HPUAanFzAsaN95eber6+BsNCcDCVJOJa3Xcf
xB1SRMWts6kMbGKwylDCUTjUygN3qfYKzRplaoRgMgmeDmPTAk+PfqfqdSjLt1OAswuASR/Dbsht
U8AHopLKM9BDckraPwyAXS7IvWqtyaRb0d9EoBRB4uk+88aqENWmgAVuyb/xJVOmPyjY93CZC60/
aOUccokPI5f0Ftp4AChjawlmah017NIbFNVFtdyuYt2qHA9Wxgq5uR2M44N7tmzkw3+WW+5PaMsd
w4FJ12RZqqLARvrG3K8V5SMps3cWteWYaV8Xlkuf7LRzJCkghzUyNOF9QVIAm7BfsTEQcAS/r5q7
/0KFbQ56R6j30hQVGM/fcCkzrm+ck89pdByerfJm4iw61mOeefrQPXBQ6dp7TNK7do4t07yRiAXn
uAv46HJ2DeLs1sHaTQJshJohxniCvVfmFO218CON7QorpVJChDeRiwaNh7Pbx3cTCm2aXbMxiJjn
smPzLxqGSLKSdJEXrUHImQHbr2kT2OR/ScVyn9U0nuNfyWFu2P7Jxtxx3A7JcosbcJpcR4JT62up
TfQnzIzr6VJHPnllpeF7EzylQMIFRjE3d3I97JVouTD4XuTv4OOSkyURyEPM3K2ChE37kIgciD/G
608q5eSDhlcSd/izjYEUoQGM5z/0Glz4gTlVgrRTFzTeGD6w27ChruAMQtlSynmeRQncFj2lzedf
fstZBBR7GP5D/2zv++yB+M3LtVXbHHucM66wwMafZix4suOJ7Vd3O4CgFLF44N/3/2DcctGj4b4Z
ptLuwB4lP09oGPkcVI+Lacqwt64to8mW2Fl645n8FsUUayXxek0YqSZJs8aDU4IrnBHozFK0NxGS
C/JEZ5+BX0qYki515gZpe6f90+SFOpTpBuInI4QSSHD4vuZnFusa0+1sxKWsrIcx+Bc5BBjQeCRV
qoQdNwpZeDTodE8a32mR/ZiuFEV/H8lK1EMhDtGfXPjEIdvp4hCHXJW6O4CTu1J8yxjDfnKRlYtY
69Goi0XKb2VYqFFU7QxLfxpY7Otq8lKglAOn49lHq78R5uRZ8g0v83Bst/1Mb9O8Ogs56BabZiAt
wNnfUcKPfstH5qRQm0tKspAy3Apa4hMI/AI0lEZNUFLodNrT0fbpBSPfyFMhYmcjghTASd/1XQNM
TAJlp4ww4KBYvWOjCiU0/CEA1Mdf/YwVw+ZlFhDAKVfDBrgDQ9vSohEjlRh9RnINlTLf5zpXvVfJ
8R4u9L1crBOlpmxdas/5+fQqGmAIT66oHemTjBNLHteL0FJCFfGchnKjHLUA0jPPqt5ge/v8Fdrn
hjBznNY/Xqolh88stPUHj9tm1ZC+tpVuqwUSn/VqaJP2IYUAJc0/gZNJFuMAaMaSj/1jwypVZv/3
zE3EwKwuTeqLE1/m+aRb9NRxnYYdyqvIaD4pHnc+W50AilYE5EOoNRIWSbvoxdMuzXW0+jDjJvdU
CmIMGxEppGvqTQoNvJ9Ib0ZfwEiHgIna0zKCPExciM03sciiD1RI3+E/mMXJs6f5jl4VL1Wt0Kol
GxEMywiy8i9e8vYm5xyE9ioujuh5P0qDscqj7VAT1ut9cdlWdLaqVYh2lcl7lLfMqlI9gZ+oQIU6
N8kkAQ9k/F0kT9/jYnj2vLgM/sRS2gq3Fw/pH+wHb96ugzyJ7a3b28PsvRE0rrH16Ew/9Gq7BH1A
1S8WG4AfCs3nn65MzbFX8E/zD/zFOpFXSTcStjDxGaGbUPu87k1n0pTyywQCUBTh4+WyL97Aoy1D
u1TBiTMPgmUO4ZKI9pC8Sccs6/igUhSxAFQURv1HyNtPdOnQCGpwaQTXJQZ4TmImlhHY4K68Iwql
GLrTCQi5JHmLDGpeTN0z02kDtHnkRvwK9u/GeXEGgx4b/UOZog7AkuZlLdi6gYdKe15nvXNYH6qp
wjdThyjNycCoN5nyDwT9cNo+V2yBZHGpEu/4SYL4CQ1UF8zk/tdUamLPjuWO4evn/irj/nsVi2uC
T3H4o60r6etcMPvggaXKG8ihx0ef4hjc91KRlF3e31rQZAdd/K5vtcM7unk/FygHr5e35b4Y8PC2
i5sjFYlDblxyZCXEcbHdguQa0s+WIML2QeYavOj3onOEzy2g3O+ElXLkeEdZXY1+wFYNKhxujhEr
Ut6KUmraAyn1mhKoJvp/gOo2dIGQsCafubLvprcgYnHQvY/X7H4b+AkEmlmWqT8CNRNRbTcEd7JX
zBrK8vCCL4JZC4IbtPU3Px4Pacy6+VCWFiEWDDP3sra8gRCKH51+qZtYomYH1gPiWgHUFclUdg8h
1ckySziHgSrHlRmRJUNT6KHOjV/w7ovNb1VvSv2RXYZxks9FzDDyBCqkqo4Q0pBWqgoqoLZ/o1Yl
RpL/sWMiAtXpXkgH1ycBIgZzH/epexzbspK3ChciHZxD4n7AzB5wrslI0S7DLAHKMCPYLX/qOWnt
A1IhfkGcGQWwZn24+Be2IvkHLSb0iny28uQZbspt8xvBTbix3k/UEPcdJm42d1ZNTSpB1sFTfzSv
9QZafAkl9aXDeIXe3AtPWdAlvk+gOHzSdeEcVP/ABAxe+WvrZAfyx6vVCWnv1TA8fWHjlR+YcQUS
2mZx9L7jpv9PW+1r7u2mPZHiQagjCAhlJ3qLDDgr2cIZST6hyODQkhO8jJ5xJT8o0d8+2fSkaGw6
j9mf4ZqgciGLPbpGAwT0VjynNeOJ+EnIX+9VTFtgFolhGDlTxcfFjBak+zYbEcHBTkY9jXAisfhe
/kHI2ji5zjwtt0/TbQ3rlH+dnJGvyDsi06DT3dLXs+zr7VpneOfATjFPpTKLCOrbJ9KwBpGY3S+n
J2oZjoKqHnPeeqhh42jjJxxjoYsFrCdtS4MnAODl1Nc70jKNvV9ckYIGyXQG87D1yjF28BIcpKT4
WZDJ0n8FDK7yN3QFqm1/WDXNDg6oJaWvc+gzF5P+Ry93azR3QdXAy6tdSCM0R85WqiT+HDFrkKTH
hDQIn2+/L++usf2NTVFPjdXay2fYhYtbqKbA+f1FqGUABTqL3NdL00+kOgjg1ZRs5efDdH8UycuS
+sZVFaHyKIJu3cKayTCVf+2kxF4sty1gdR6G/ZfM/CRle3YKeYVbhev/5IQNA+t0ybfUyo+y1C8q
qlMFSf6pa81c8n3go3lPpwqnI94eEQ9PHGJ+HXQwxELb+yiacWXebaU9uJB41GktPzvPkTf6cyA7
S2JgnFV2yF2c06xWeDHQzOg/omMl4/tFHpQaV4UJIdv1eURrc/+bAE4g5MDMV+5zpolFfWR6efFX
1kulbcKmQzIsViRiNtyR2NWIpuMj1xnaPag5nwlkARWyzV3SbDcuy6j4R/Z+izYWgjHXPyyw+Nrt
A9PrLgjWzmt8dH+IfpCSAd47WpqdswmBh8/AzGq0dvgKoyh49/Rrr13sSwBvXFQCqUhg+NmqyqoF
0+73EbRiphX7/sRwdudVluJ8WfUCctA6NYIDLCSxL+Nsw2+xGNXy74t1z5AXXweOkI7mxpfsMWAM
Q2Ttum7/KZXuoRF3/4C07dU8KgQgg0Hd1WmexQ75pn5bG3G3jx3NA//MAScCpEeJBCRaiP6FP1C0
aeOClGN+97p7hSftkOlQLuYpwJtg9OOqaWewahEIN+rYKC8HXfPEosL2oYP3WLYilk8UdJ38fQnS
Vpl4RAhxR4y540rguJG+ewiZE/IR8Ayt/H2j5ibvgWhDZluUFuojUIMvGI/hzo3nBzdHDRe2frKR
5bPKuAYsvrp8UHkZOxNuGO136Wqhz6J/VvmVOLJFfkkuVPBUkNvga3s3uoLu452QRhsSebV/BaH/
7//pfhXlTiEOHX0F+3cfFHRP+ecSJHblgPf97y8N41QE0e8Cn1aIHH6sos5GuxPytl43EoviXb/7
EQxmmZ+oErNIbaSKILE7AERDcqncZJNNn3jbbCoJRBoiHP1yaNU3fMEZ5kaSZsHXqoZ0mFxSVMvj
gpAYr814PaHVHR6p5BKGqZEtKGGWBNf25E9EmRcQMsF4Jov7p3MEufeu6hD2iIF+ih8nCFMjmJXd
h4tKZ9M5x/kzwyYOIhgQ5DEcsC98wWvVX3EElzodfcceTBbkUncnWPFMHqC2kZ/NwrwTjKXohOiy
ea6QiuprnjfGoV73O4FO1xs512wTIFxBuQf44DUDceQUgXy6vDyilbalrvGKjbEtqUkpSmXZcX7c
JuaUwa2/QE5o5tG23KdhMuVJcw6+FQ2ucmBV+HcxpFlF2+MCJGVPUJqcrX4EFG9uZEfuEAOqQQdD
CD4eQ4FCspdPLWR8FCMCob4EwtAZK5T7VL5DAHTcz4Ez2EHvP4eqyXOp4EzFwJxnZrQ3X9sKBHyn
VhHUcPr9QexPu6Y9WOJE+rQ28WwlaTwS74WSVl4zcy8JzytVV195u23f7lPXK607diWz4QlA0pbX
OD4iEH5uhIjRLmjpIWcLvHRLQQfjoDDh1154iuBDHfu9vIbiekhPu165/17fU0C0NvIuWryOC+x/
h/aOKP0doSsqlH9HopjqD415kCjxds68cmPXPkGS/YSzA7wc7e071S2ddZuUcLYacnmoRstuxS6K
Xmsx3R3AM2uPIgXhwWKFm926DPt8cpkXgipIEl+s39y9cT6R2keYDM7r84l4kHG6CaONm+XStMMW
OdcDtcQW7nUFeeOUJ1Cnp3UWv5tQeEKTrPFnqEWFb56UJPGq6odf9b7R83kvrOMZG7GyoxvydLak
qPfbpDTEhl63bcrWtvN9dj1fTPoApg8NbszWIIHKEwreiZD94NRwwUDBTah/nIkCdxRyb0/eEGXS
O1x3ktz5nUtoGAaCWx6cXbFfXfC3o4+MlqtfrAZ4/8mK6VE+XpklVsdr185FUs44rPaiiO9UdgB1
sLvEX1H+bQ7lJPhWOdxj/SW7KJUaQ1spXoB7xsm0MLQM57w14XPnSVvQFLgQjA8ZvTE+OWdLXkzU
rKj/Ddi9on6PKryop8H2X3rgP75BEafdSTlIWzG06qn8u7VDMSmLb6vkuviAu8HUBX8YTidj9Zhi
9Ucz2A3hn2a1fn1bNsDq1ZbWYo5mFsAd8dpVkrn89HCoh8qiOeBC91xAU4RXFF8MLgT03bpkz7Rs
Amh0RuTHhwJSDiTFoGa32KGpeNZQJJBMpKvxSxx9jnS69QXvxGbYpRYIG3c9YxVWlmW/tr93+gMi
rIp9KWYbdMI+iO8dTqpNplqhdNdEhxfCL0tH7007rWw/Cz0P5SU3HyufZ+bH9/oy/F31mJs87AOA
dvkMS9tHsIrIlDV0L0gvyjZ9mZzHxQPRDE/b1W6cY8xDFYDHeiI7j2wIwnQXdZlS2ao3Isg9gEWn
s5eGS13xFfD6cKSwaovOHijNfEin9LanEV8lZZ8y2uz7BM1UH6JqhT2Sw7O+MdEB7BMD+rbX6Ks3
RoMrL3F0BUExO24XImPrRQk5bpaH3SWJ1l3UTCcjGESOxdrDKpYnxUn217slmVMI8ol4BpAW3KAj
3uXEN+/o7nkaX23BDRBKMZexnBLB8TNFigwOuLqntOpvHJ4gumyp8Km3P+HeId2wLLGGDSkshZRb
hsG4Pj2GqhNsSbdM/JFLv29hwXZxF1I/4h4i42jvRWX9KopiNuvtSjRl40845Cuna01TzZ/JlQU0
fl2IDnctfH2tUwvxopt9VDDn2nsXca3ginD9FgzP57XZoPmdZmW5tENxkz1rxgx1FdBtHM596mz/
DT5NBQ8c4ZRqs6/DA/+a7znemVfjOqePSKzH1afROjb6e8IfvBeEtKaq5tER7n93JfCV8jdj2X5E
w9sFhk0UbPsb9vhcAeLM5NAl6PJXD6mOg09GLwrVeulbbq4KkbxX/uCkSbJ8aNb+rCV6eBxlVfgb
bDdQoYOuWpaVUQZJLX1dUrI8elyg6qGB7kVizN0p8t52jajxX5OYQndwXsAw3YyDtqVmDKp0VUX5
e8tJ0OOFjbUc2CiFGJjnQDD6coL91DRu/Y8MmbUm+8U9BCFVQZaiDF7hO+Kiy30IqLx/hNuaoFN0
gt18XxKG4dTEa8O1jEqE2i7kuCZkq7r00u1/dQ9RoNXwzzCi6UW1nBpKpdDGCUnbSFq4Rh/e+34C
G/Z1ZwFMovYQRgRVBwol1JXUAT/Mm6dwFNKXatqG2bjMgpxrKFvrRmXdc0k3G6kTR0VahGevkByu
lUf8BFhp5SFV3vDN/Fpq4OMFnmMmDAptu7ww7Y/cm9KZniiOIprswhyV/Qy+/XKUtXhjD/pSTyHS
SpE9kqR1bKW1i3WSLkCt5QYVW/LNyy4Tkn3fmrR8MPvXC2CQb28fgCJGU7gbSzsULTmBzuOPhsxE
rO6TLc29PrUIrAvB3Og7jsXFAMkE4pLzu/tE7JCPnkoVV8THf8F72xHAoPPksnwlJ/z2GprE19O/
xNb7MnJz3jsJcUtiDc1WrztXSyG8AcYlbbPnyu2pQJ6pfpNCgyz9NGUlT8O3NKccGcn8pkdMpL5L
A7zYKVi+w3k3Z9E21aJXe4dwfzkU1pgYxdiH4juymuFTxD4MbFEPLpQsn6vu/QiqvTdAryGfl8df
od1NGq1u0z4WyW/ImLBRLdJRulD1X4WgzKdloWRIzknqXnaPWc9WA0AfbowxNzHh6UFY12o32fpc
7gckvNBYzYOS7moxB+bu+iuCbPqeTNKCL7qCtZ1yMDGKmTf+EBFg5L5DzrdyFuirJb+lv3szQ6jP
1uCQFxP3wFipMgvakmACRIF2v1F8tDa+S27LFNwxpxfY2Cw76IeICJhrILs3ZYFcBoOfkLO4i3E2
uYIhXDvV3zkxYYoqj24h3Wqi0R+qHC+HaKaK/RFkur5hFbF1gtIravO/cTmqUBHrt26j3JY/84AY
uURYBp8NLCoaJbjUsSfTQ9zGC4WPloUVAj0z72RO8u0GbwSbmWhMgJjuL+w0J9zpdBeQ81Ubm6wD
j4XMJAS9Kj1m55IcvwWB/G4IobCQtfjfBCoADtQEUsQKjhfIxMQ8CJtLA0DwOD3kU3ZY06eKdF3C
aZOcUdZI9GkjFSGWipv/g3hoXZPMTnif5/AZm48LMVgtTFawEpHoqP6yhxZJGHhT1E5HmoDFAGOv
axoNV9/ROrv0YnSj2CgmxTOtZJLkHxEZIeoDJ9RfU9V1KqxfphF+b6PLm3EJpOG+foGXEvkwhEwo
2b28BeEKY+LCV8w1+5ffan+QrvphKeXGyT9v1EUlFCvmL3vPOuhB+Pp9J+tnc/1WzdzOIlIJ2Bf7
8S47MJrOo+nn554/Jam17Mqzy6MeHdEkp5+iFrGNrjZMc5a0F7F6q2GJ7KpmaeiTQPSyql/Ea7nx
Gh/sKmf6oQVM3vhNbo24BUyZzII5TA+4nzX4015neFkbf68bzPqOfxFMqg+r5Z2b9tde0BMhUBzm
XjTB5m4D7jPUbLldDnRt3uh+sy45we0aqSXxphLSETWGqY5VchvUdhi12Y/FW4VZSf1XNDL0ySTv
x021Ju0Dxf+7KWMgW3AZyq1iDlx5+/WETp/CkjYQGUzc1Z5FtA9aCz6NWjfDWm4s0ct2GJzgkztx
sb/3vhRGXe8IgcbqWl7RKj1SXt/G+Ha2o1T4cn4QT0RNkaQRxdVa6w/fvSWUW9SKieIEeuNsFxdn
f4I2I5123/pc++M3sN8FUdYdevyheZqWwGxh06z0VCB2EvGeeE0CAlq270CEYHHT4ZDgL/vTPEUz
xIwho6cCfmzpOYIUlYGBxj9/utlWHZrzUwv4AZf6bjlP2lsqUK7RIxHvKQ2D/y6gHmqmjSjeisdA
gX1CGJzdvrzDkkkLFpPrJAXdWEG/84DUsePy0q8w9/oaErEvPrjQZbzIEhHkxHEXq72HN0MqtESM
qR3YzbkDsrbA5A4Mbt3UROClLJr8pa3Z+MAxWgv5bLcGXvfSyI3YVkxMJgPd0CGa0tnjJSX3hEKA
PcEFzTYKGvR/q6EGEj5RQetBenaozoi0n1nPX8k9a0QdWOVXEAvRLA/6x4adndQECPtxP28sxIBl
B1iphs90zEm6RczWf4fXROspa7QP/xnFyS0/MCEwytAph18ZgKwS1UOUq9BbX2K7DP5fc3MmXTEh
tKwD+lwpUX5EcioM7SRBsnjVueEpoIdKo8hODbGYP11/XbYlnnMUOcoB4A3iyNU5bp2JJ2e8GI4h
aLfpyyuG1AXxag/GPG4W86sBxXUcGwR4p4pA/SzF5F/QTJra/wmiFMVSWluQuA4nVOHR7L+lRlkZ
ArX5Z8pvDBHxhizXrL4G/FA5Xb5a5HVgsDsqkVve1WXiRcO3Tfca8kRDisKYsQP+qWhqGesNLt3i
dFVBmSPljkxirXyJeJAWd3opYQhikC6wpq7Ldm5rOgBU8FafL+krKyCGZFC7ZhbbFUQPGUcldLCP
1jnTzSatesF6ko1t6/XyuIOJJ5YmkIpp+JxTz333Gu232B9xK9jiC2fBSfv5HMPo1mze6OwVC0Tt
vTl7mlCHPvXb/wrH5310V7iolLlyMxXsCYfCqlVfgFVHOqipxj7HxuxnjTR9l91TqkaTUZ3AO8U9
NEw+WLNr8A+8enk9X8XgRoelTeZUA0R3Ool2Nznnyeysmzrlklb5Mx2hPtwm3p2rm+D59a7a4eEH
hCwxRPGj7N6NFhUckofBgqyrYqY2zS5D1hbZz9S5N6Y5ivIZFLllnEysx5CcBk9sVxJFSDXFdaeg
dFLBJHZFlG4S3Y06Sc6yqQKf5/X+ccOkhwdcnB9tuMeB2nLrxbIPuOg7n2JK8AHmiWomNOzGf9yF
38WQ/Ov0K6aG2lnB5JRKXJwvZNh1fEt13NzJ3y7SL8LnT355rF56meDpp5uw90qydWp13OVfkyzR
FnJvP6kfPbhajvkEs1MvLxZnbsYn3Z7K6+UTH1pnzFf/CVdNkqAKCSSJDtwYMlaneU4jjmnm5/Lg
kgzNfx7Q9dzQfm3YLI+6b1B9/dT7wtWe81vYcpmZSj/b7DKQPUeXB+g4+GWL0qPIpOh0EEYzrID4
d+NBCe45fw0iTiIav680NVWBrWUekgPXbUsQasHeN9w4ndF+PElAN9LbzKsdP1/wfUT1v8zTlJUq
zM2B4pDVzFG6Qvx15cAy91c3Asz5ePXoRzCDI9UYDXSLIFioRNjpDR0g/6sJs8uLQrX1HCS2zf0O
EIbnXll70atzp9Yy1bKfFZTa2IxIqx3dm7fCibupqRp9RJOlA7sV/cLSPrvOW5p0fn6H1OG2+KSY
77zYANXQbTw+lDSqS0iGLU6DCe681OV1sPGYqFUwKlRdzlHXkRJBqOhqQhXzg76iDAJRA4iCzWaq
jUELDHEUrIinNIi4Ris6Gq11yS8wQeMUYf9v8CET2vDjPUFbAZ22mDXoJBTM0ReRbBzylycTsRP9
Yd6vv/2T6FORMz7zVvH69GHCK4vTeQHB50hjjnWAiiFUEkSgnjKKrWYWJQD9ElGud7sGzyviaOfU
wz2tv03pyEZPtrWv6vIFOvP9jWZPXlfLfzo3fgMLPfzhCj+tLkfX5nwIwDFSR84P7Wn0tHJvomEU
x0Me7aUiRXY8SdywcgcdyrCg5bHhv/OPJBN1Vo1FokL5+yWq1tQWPaGeqzxOIgfTwDi3L/ZMHkKO
dT6lrH7ltRIZkh0eD5xfiys+UWIEBLR+jrRIJtHISdmMYl5P/OUBKqf5vvNIvG6IJwXvqC5VvzMz
tJJNn0O1DY2nh4lDvMyfMBSkXULiy4hGE87bqj3rz8NLmAveyqk2BE9Pj1GuM6RcwC6GeuZU+JOz
YVrNNv8boHzZVdIeSOdsHG3Wsepu53/qOxWwkztFNvO9UfkoYov/9Yi4XDp2YySiosTJ+MlzRM2p
hXhS576AUvd2eiKLORabHjL4vmra1rF5GpXHGeK8vDle6kkCPTXcDRVZy3NRcynCezi2PhWhDeCp
/o73pTDnCi8RcDZXr4/OKvEZXtnrhnL3gEwCiiqImYKGvAqp32dzOn5CiM8rgAfeUzNTvSJe72cn
FgXI2qH2QxDe/CYghu3Vb+fX3wJg10QTXwpqSi9cl0MgK6Eapk4afRc/n11L49DesAkXUVqeOsBv
AICJhI3UHYNtoj3WgVqoYCn6jrL2umyo6OJJ1wEivnYANqWS8likTemzZLITxye3EgaCtQaAu+be
BhC9hVa4N3c/MW7xNNOdPDdFyyQxmaN5OVQywECfHnECY/DL/n1x4yfXZhned6DnK39T1aXkweSO
SXRjsaxU4o74+PVHlSL+yoaK5H/0GTMllNTTur2oaYXs0r5npRUc15EXdtvwoQbSB84gAzpuyrY+
aiSHOagg9p0V+UYTVQ6Rq3NR1Ush6zF3K+IyqhfG9B32+9BZLq3sjmlSROAFCAfY9LfK4zgpE4U6
ZcABGByPt97YKjlzJgsXRJn2rE0R1UT/yVVBj29CgjG3f4l6y9eSM60ET5MsAku6R9y3wH4uGAhU
9gDLut1CPfREWX9YDw2BjSRvtobO0XIXCHOlfmGl/e67kVXqHOqGnliTzLP5WCFcYRNbn8gV+B30
P6HTO5930T7A+pKs1u3M//dxw0q7q1qPhKW2yB1jGvUZaPlxdqr7TMAZQw8YsH/o4h0uvuImYJR1
/F5RsQOL34+UnmKbqh1Wabav4XrU2HrW2PSTbWEAzuHBUaq/msy1gEutZkTY8f0rc+ICWQsj2CHl
cdmcqheCYIfNzBKi03V2ks/Y3l/AUTrql9s4aX/fbBLeZ9g80jJQ5GJDhccPgi6MFD0M/XQmS5gU
9T29SBGwIb/os7hiiZ4BUcWxtkk4JecLrVvd2EMYq+4IwYNCxSDp1N/96q4GnCWMk/JaMqde3vRm
v4guUzos3dCOFwVG1TRIzLxGRJZ+mUdJ58G0Pbt3QyiyJC2j1cv2aHmbJpgLSUni0+WIA421gKaD
mCoWSMUtgzRgFHZuC8QvLhTyoQde0QAYNM4rLEwcvBjReouVCwiAo03/e9qqKYNGnaF0ECMhF2Kn
Dv3nUQyH9uPRW5D0n25kMT1whldiEp6i2QWOF8oiJa8bhPfAlThoCXIgc/ZuX3Fv7u2Wn+JR7z2I
m6Q2jhynv2MEl2FqJmdj013CNOjtlDBeE4RTNMhkWT3qNc7ruFsi11KLfiorAThboIyNloIEaHGN
vRP6mF9y2FWFP1dK0FhVSnF+3r3WNFal7vcHA0TzDOuIhglvcreUlRPp3siOmMeVmpwyeaf+Hlml
aVYvLaDXmDeNQs4PGlMTCdwH65vnA/leLCScX02BTVGz9Cfpn7CsJpLqkaGnsYS6tBrWnOpbluWF
ugWxjLRksPBi0LFtXeGkIbgZ8iyh97MKt0MlIe6L+iGlRutMHG/TBSMomersKfzJQK4de/wFHTGj
W80kcRQ6cJHJZmXGs6/vTd47io8hBRgcBx1IL9BGbyIlzJyOpzMV9uE/a1VpuZc6m5tjZj1sbtYc
PWMT6BK1n6nMikFq+G3Y8Ca35PV//6aq6ARxYcMua5UyLQifM8l0vPFIkfdz6DKwhziXiKxqnK6y
okKBOLXXvgBeffGz9Tg6YHg6N1RDnf/8KRILI70JshvH/1lNXiXDful7ybTyUE7uqaaskWToMaas
fc5QkdFMbhu523wWdotEODStIAyTLvz0j6M4lvopBbC9AqfNFMYGEHX9bNhsowl26BsXoGOycF6C
urm/0KEBr0wo/5MXcFwDSIN6fWpR9FzoGwOHKWB0h7re1pmsfWh4DUq9me7JCbTcT2JAmt6jwhbQ
m3zLoMwdtCzC/jBD4/yKjQVC7WuPgqDX4lQKHmkTaRfBYxPWW8cTO9qNkw5GXgrm8s/gPtQFtDuI
uIeBR6CKQW+7DLM+qMHCks4pdenjQ/hZsrhsH/V8oh1Tz6YdppFIXQFkwjD7oh3gCEmADw3nPi/X
UtJ4db5q9A/dHf/yI7VgGev4D1JSTKl5u+TVbQfyWnu3hj3UDpFCvlugzsxpPV91TJRqAnv1kKyW
78UD/VNkb7g4WEmxwsexLYOs1BxphABj6tei0+fcIsxWdVU7I838I3OItqtTRtD5n6QsI4fupQUE
E1WT37VnYy5OFNjaiMV5Hcbjajz2+7YNjwJjMkeEkTclDXVNx9F4XVGGqufeBFq0CzhjqqzM1Rcw
hiNwzx1ZkIIONdpYxcU8VXAJYK4ro/xPyUYL5YX3ISfj6hZOgVvcX/7QQEqfG6DheYUx7XMIkC8P
Sd2At0TmSnUVXVoLsM8bhg+NeXvuqY0WUe1PJz/XK6OOnvBnJK0ME22mB/2FpKeu+5BklTSqBY4/
q/CgkRkA75KxLcdQls2xkUKLRXgohnd5GQABPsmpKqpNw1o92eF1WQf2xph15udC++GYElpc0QZV
P2DzCcE/86+UZ/MDd2PVgHkFyGSYZb5XDBzqkw8JsRWwluMG8ynkIi78ruujMJ/fub6F25k2MvV1
YJJRGpt+FFzPM0FXHhZnviVdgzAekV1dEDAeCutVD5o+ARBfzxEqiqyst3uEX5VzTfyUgnEFZ1OS
/25iyTgLs2WeK2pZfOw9NvvepIAcE5/a1tcS2Ogc2lOgaz6XXcySkVmMgK41RJ/47xMwa/NWWRRy
qO57XH/n41H2Ipm1kcNeW1slSth3UhXtUnTTJnvwLrRbilDSNMq8yUtvJpZWPVh5COSbaMBWV2p0
0uLps0wVqqFO84RWNG9g3BQSftSC/F+sUrrNruG2U+oLQImjyqLO3DODmVVs1w+gNvrzhm61oLUS
Arnk7ZxR+79UOV6wtJRcIcwl5pnfDCQw6g4pdHJoRi5ZaTGblM+b4xMLRhH9+4/Up1Kd0n1ibQ85
PdXQrpRALqAzZhWXuU9opWg8YdVR2ZsXf2A1nHdlmg11SgMvFLiYWYYi8jXpd1UeIRfpLOT/mVmf
a3aMlrwJm5nK3tKSAsU+3lRrfFq8k7WK2jjG+mEV9w2WQwhwubJcTBlgz9PXwjSGHK6XAqI5AdC/
0GqWf0ZSRcMCghjQ6VyySquh1tvoSXryoDPkH5uxo5CexZHlhsCJ4AFYrcHVRJqDqSYL6fSUyCGF
xWz0oQeY0AWKrB0cCf93vCopFczMZJikhcDIfwNzGs6z0hRpj/fQ9mf2KTLDgGu6anezEnfh2QKi
81I1k4MGAw+BmBGRsdlEkYQmroBnuaI2B3hOFAnXDwlHK42G9NGu4WwSZiwhjEZJc7o/DIwFvUuY
8oQmLD0mxmG489m6Q3XOYBN07jzMcZWGWP3Zv51fOwsnYrrHlRLrtVnpPQ8G2STAi6kCnyHErdt1
XGoqmGvpD9//k20IimA0YQ0Zi5bn/g6TLh7i0sZiWTtlnz9mD21gnqQtO3Lt2iucXLeev6VUAY4m
bLVc/iRmKE8c3r1tAPHiGaVJ0tywkAHZ0Vh2WIpsPfwVF/XUsqJQFTgiXlY2KzX5MY3QN+n3aVfN
1Z+17ewXnPkiSnj1IjygBnm8whcLrjw0EvJuf6u4kO2sSfFX4lWVq0cvCZ22PEI+7M0FbqcdCpje
+WbXoBYWE+6HYkt6YC+IkLZ5SmOzBhGbEM0IwIt9LSFygQOmbQq2aFVdhzTyI9Hbeu8DuF1HVkWc
NER3inVXibp6WGHuBTFCsmsHrkfXG5gTqElk4oXewD95K85mafYrmdURjL5ymzXQw1G/ed3xdp1t
aBuygdvVBG/e1FGNtVVHfgGhAO2V+u1mGNON7Wh/cMUAAUUfH8NIrtoOvOCgtVtpwFf40Elzg4iW
YoXX7J854jJthJ6JiajU82oBXZXmfBBQTLfZAfgM3cvc/XKOpNy+3TIVLHYSOuxzo5deHxz47rxc
8AWPYeihw1IAmJetqtdbGK9cqgmtp+722UktuLLXYOklibiC5wwGlVkaYXcX38TiEXtg1Qj8ZwFv
zdQF+eyQX5nsIkwhxpuKsZ9wQ9qwyCTYbmHUcNq9JB1jWNZXqVQeYCr23bgN9dfuVCWCOCIsQi78
X3saR9Ic1VLMjLZ31pX2Qh+elJ+AN4udhmO5OA7J8Op8fvjg+G9E09hQS+VG2Miv9VmKcTJErmig
2jupSq2Zh9DNUV8JvUYgjgswuP43/3/aRzS14kgC9Pfx3C+oz8Z/xw/5YU3sDT+TtMgt04opVKa3
BCD6WS2a/raFFTRUhSj8zFjCPOSpKXoXQJymxgNgb431thysO5AQrQ92QcB+jlneSkpaBBb/P08r
eIPCEGm5LsPk+BKCHSRLtEZto9oe3FGmIIQBtRuCPwG1Ol5Ykc/FIDOhCBpcVMkLdcbcpaDgwit1
g/xhB5rURh5YAAOv/HedDlzKPNmaQ6CuSCJrWHGoBK3tmc5hDvpGECIZETwh84ETWdsbDbhhYLWe
7iWulcqdbJfpJYyCslBRyOIc7+8b2k1b5mITO32Lq3tY87Y15BBliqJuqnJchudW6zAFrK792u1J
BO4iG0oelH6nFiwcukafR200laQV+zavA+rYPa3cnB5Y3kSwJFHVcBjN0vjfr8NaPGjAx8VQJ+X5
QUgc4UtJu3Y4ICSgbd7+7lab6HpaCUlyOgcNwawMzCh9Ni8l/Xkta8xD3Rzf5c3ZOLoV5+hqOBnX
7vamn7VMAzUGZA9KfOTb330ihfb1dT0GNpUSvbJnvfr2p/KdYpYVudfJApyLe5bbPd1V6dRBhkE6
NvYnAR/vLmE32WDSDJqXoH0cOQldhNgYWYF0hMfzn3g7WKEAd1jEuFFfU15YQeauDmhxk7BwvIf6
/QGGwubNzxXeh2KVj3aksnbzPrBtc4LMbszaqjfrG7ci45+ethxV04JJbPdWPAbg+k5A0syWNkLK
VciYxX5vkcCSYG9fNz3CL8r8ifQQZvIb91uFmK3H+G3QPoRIvmyeOGOy7coJm2eQFvSdBDIb5uWN
Hg8Q8DkkX0ReZy/bkzR9ffzhoGwgSMr7lWRbhfJqGRfNVAuZbbkJnuXG7unv07nLySbR3QIK3rYL
Zvlv+ZjWyE/gyHGWFvIm5aTaHKJKONSQbPxF96tB80KslKt25u8WrczuomggrTe9bnu6dIWEHHRm
cEB6VTMKmO8gIIdU4boW0yu5WEKtOjQuRXI1TyoBtd1zwDrT3rf/XPgJDhBSwoVBPEH7U/OwWmjb
g5aPcONk8fl/JjHP29sVTyYU0W4YIPGvR3yhhx6wJj0T+icYTKEt+Zym+V+dXMHgvuAoiOsDmg2l
j6l1ugyDlrvC/FFGVld8WsWwAlLYlFjcenhIjPdo7xc/wXp1yYROaM8Vv8pm8nJ85S4SM/zerP38
fUzbU1CuoA4CHjLc9SD9zN9UP5WoTxpqkPYyJEN1cBk5gvA31Mkx5JQV3Iio9uudNsGcuhxIgFd7
ciqpq9KiqLUP1zixn6c+/3x6L261prtEQ+K76UQ3rxv3aAJ0gNaxx95MJORthwAUAuPKMca/xy/6
KvEs2L+ok73gLz1kmMp6nvYhOdvfIXCMOowsgWewhNpa1Dy+IzTZRbSKiS+j8fOSUfGQEMFDKqQq
rTcInyHqChw4+2hbiRLrmMmr7mZ4WUXHj7R6p0Q9kfR+QK0i4olYdq1C5xBMBGOIp6BzVeGLxKfZ
mkqNrZGzukg18Hz1DIszvzW1zwHP2gPKpT9NC0GKisKTqXQdcAFt1YQfuXToje41+LkbOf9PDUny
Gi8TMx+eF71byPhpRgX166+EsxT6j5XsqGLTcqYaD958xAlRz5uYGFeU/nISct2xTS4j+aMSN68s
98Qn6D52d2nE8ukDQERmlC/2fdzElvftFn+k7t+KWTV0n4BiXdOP40ESLH+Z4GTPO7xjPQtSkJ7G
lESvjW4kOtHJOWsD6OoFe/hMt/PxXQ55+yUJxuhW+gsgCHTdXENvwCwfycTBTCkI9Rehcnw3JaSF
StAQDYTVpcg6HS6Q7jfBmtLWFF95rpOntLFLsNfPZ4ioNWYrzKOdX/5fufwerJVqvpvLP9zW/mQ5
Y2zpFoiXtj4m5Hee4/G2Vh0kzbtpoNVFfkFWnONP5zxNC6eB+C9Wf7yb0pm+SbGMFDeCYl02huRq
ThafViM4bRF2MDpIwZlOYsQGgJ0S86dYCOC4OO3T2vkLan2O3JCPjJbAPNwiX5kAc9ESv1pyapnv
2nHXNWDHPPWXA6e2tAbjgyGcHzBDBa2A2Pka5OPvG5rf4SjBCMbUex7B02oEzGpRIFFLIrSR124T
eeNox5xKA6m4IP2E2YRiDm+xw89UeAKxUury21Br2DNUrV5s7UTOdw4EhJBRjRN+gRb3GKWFmKrX
sarMD6CBZ0/pQWUV04096KfRfi0hPEQlVmLIIE/gxYn/AOtfzGYOV3rSjQ5JtxEKsJ/5j4ALTNZH
4Aln5YyptIRgykXBB8qV0mtAqLV8VvyVQAKpsGquDBnz7hsKu+t2Cvdz4nFe8F9T0x/xBnU6ETvi
1xVjbqVkMzfY1M/V1Hp+tRX93RsCSY2bFTypGFy5+sD1MF+FUN7pgQ+5IdVL+TF6To0Gd+6bhraB
VxBLzU+M+Q/P53t3cuEgKFTsUmJswJElrDrLgtKQRP1Ey5fRKF5aydbN/JvIPa5p3BdhYvblZlav
guMQJpFvbvyjxx1Ov8j7f7oAxDI/TmiWUWLPzUd8fsE8Lp8Awq0J96He1vWN7XGjCd4s04+g0fnB
xp2YC74O0PtpCQM5LlBgUyxZ0a/gqCAZACf9DN7IUSafFeinAV3CkwctsNIaah5IZ/uLB6RXLVhq
wNTQG3dL8v+mTFj4X+pyj4tSXakm5OR1+yt+33gZOsKV5m72nfvnSfW0T71mLRSxEIICl/SJW7Q1
57v1imbHYZfAVXUfYPlpliXNcyxbxV4dlb6+DkpoqtayqHBZ6e+n8Q6xvoe0L67GigaeE9WJYthV
l9F4YlMYg/JZdA9OpUjaNdyXO+DY9h4Trs7T/xTFV6ZKYpz+oai1FFDx06HSw4yjIxtCR5NrUOZN
PkGx+tYvGrJPBuGjVdVNol14kjX868D8keUh+yhzedhs7Q95ycNyQHgUhbKrlj99MXpeb6CP4zHW
W3rw9c3MqoZp53zsdiQKXbM0aIwWFeUwEIGnCEn2YLJC8as9+YGv+eC0npPjH7VQBwtygWoT9ghL
tzah2/kjSEutCMy/jHltbJduOGDkOnBb+MH0RF0zmwo/EOMC/43wHKjM1vJSGgBpQm4wOoACdtVq
6dLmG7YU6mn4JI+bZhfIspa+L2qFHEyIliiGXEuVelgdCor+n4o6YMCxuMG1twvNQk+f1CIfZ64y
OTVDG7fhtlZS5cl6pGt6Xc4kG9suqA4IZvUP4LUrWUdlbKUEk19C6By6LOcraGWg/kbTKuHYsC+k
6WL1zAJnI0D7INyGwWAI1pd1hfFbze6RBVe3/O7WxIoWtdtnkHvE7SanGxIk4l0Afjy5jJTSgwA0
7A0BhGYpD0+I7KvDE38yX+RKtEnxJhdTeDgsvlu52i+saOhYI335xZz0m1MhjXF2Q9vDc2/Hpa9M
dypjKpNztQ/Ax6Wt+8CTj1DE3KgRfq1UpIM04nUjCmp6jMq3qZhZR/l9h9Bjd2ZcyUZckwAwaFg6
vxN1zip8LAIjvAMwQUHbda21JIOe224by+bJC0IYMk2dmSvpGKESNxudR3XtUe24fXGbNNHsvEWt
6bkTW5ShzcHX2tXeGZcuRBVWtwYu2kVs7alkdHG2+9usvniLy7+0kNedhs658obAkuF675Myqtgh
ZeqF/Gz8MjY9D4v8T01lPxpfa50y1hngmSKaEh1H35HIzxyl9Lz6Oc1v81aGW5VvL7Ijla/GV/wI
Vs1dKMvF9QWYFuS2DwJ+aXGnEKH0+JssNZZP8k9dj5ss8yjFDNfoYR3RiwixcVOiXLMOpy91xIcK
uw6x27NTCV71oCnXdUJ+xyI/qXGPfz4c5uGrHjKo7SKXuNbUsJWs18JKBEYrKOyPdjEqA6wvSX0I
NI59brdpiT8h8PuAVusTsu5huRADuDWur+sahZ+28D0YCY9pAB36oY37WzkZuW9f3NAGWpkyIEJz
Zf7EufDHRgY88KAp+092JRaeKbYApPuRKj4kcIF19dehXeMVyZrYhehrGO4bIL2XOlgxrKyZ1RjP
NbOK8p9C+lQj74I8WvMdy4ZlzoBe2tjgi8I0PqY+q7nacl+pydAippQK/HORabs+xdpqbk0ljkDf
a/esYuNI9u7OkzPcXoNnjO/SDT1Nt4AXT45i4HlA5UfmWSMhpL8TzPfGY6V+Gay80XvildPdYdtn
mLjilnDx51wSogIh6BFU00g0E1aAZ9oMTY4QoB8LePl7bmIj/Ok/jU7Syg9DXjix3xFkUa7SOnlV
U8IQ+V48Ue1PlsM2oRhNl21XUB8kGhbUVGlFqc7vwfPNFwb/grVTMYaUF6FC1p3Fm4M8KcaZOSK/
r1mWrgyfePuicd2b5RJMWOrCsgO5w6Tqpnmf8Efc57Dg3IZq4Kjbu1JdoVA7Ha30D0TmBYA6xIhH
BMjmxpVAlEZsPLRajl9P2+hQyslNoH+5friWmIaEgiaE9bln7LsBIyXJeaCfbsglOEDfpRcc9mbA
jaXzFm7eAz19s7j/lJ4zjekvGGW9Gio5dGznukxni2Ok9ihoG1kL20uGWPCuQzenYXWX3IB+vzhE
muK322vUB5U15n29TlVwvM64RW/uWK9Wa75+7jXldiFyk8Qr0WJ6HN+RCpKDLWuueSuGjyOvTmbL
D6RQoud4PaTEoOeSmUwRAvhwrgC1wj2vlmGkRIa55IXc2nki9tKF/VpNtVBdjwOFdk9NPP4O9MG1
41kMKvSrgTp48hca8udfEQHVccy1Jnk+Qf3nDyglHmm/X5FbmLUHfZyArcO2sIUEXXmCdtsyvfZy
b6fE8zBCwcWA9P8LGw7I9SH7gdzxQOZEAhlMZDVjepvOXFaTIohd6Hk0libUQ4PXpAcN49g0luEk
a5KGpZs+Ip2GJTedjjxjmDmnzOmETvn6xp7uPXmcTaIzUKV4RdWIq6yYklKmzkBlJgOQoIQBEVV8
B4IUGvBdqhMof1FC7ZbEtfGR1E+n/ipIUoPRHtuYN/xhqc7WvTXTq9qaIifL+XA9A4JChsOswvBA
CUrBxrKDx+sCzgBFVH+qZcKHIsN3iHElDbn4lEQn02UDp5Qdjc9QofJHUY1qN1Giys0HjVNP/nrL
4iKw9/eemoYILDZ/VrBnYqiZ+Rs0WOOboihH70ldMzcO6DSQHSuXigAfomhwtUyyQfh3l8aIhSK7
EcV56nl7Y0CBiJ/6CVUZ208ouJ4+MaxaoZXfx2VXnp206jLVy0vxrQLN5Ezoxb9t4jUuUz05fl0V
E5mlFlCq5rFFWL4uopGbnDjf9r1VrwOuW08nyCzpu0V1XsG4hCTmpwh3EqKZ2WiReX43FQSm77Yw
RH5VfhBwLL5ZiJK2WeBbaYc4/KBwSswMLJQmRZoj58aO10uNeCSga1+mP+Mjb6Gd1JFbAjtZlV2i
NI4VJtHBQUFjWIa5vlFhfta04wg58T8uufL/c74ThNRZquFrR3TuL1IE90RE9i4HFw005hCRpnhE
P/4wWQroUvB2hhSAuAPxxRBvROPvOnUNZ7yqmDGX1G6wd2NshNVewf+HWPl0EknFvOcmYTKGjMH7
dittkmqvyApVU4UoRjPHE0Ido2FucsBuiMrioxUOnmfNMBlrP7eCfRhRCosIiJ3A3Y5hRUyRPEDS
UU8PEiAPCTmi81rqcI/nCyauAHNlHsBKk5nD1YC/brZRqtJcp1gpTUj2E9iZtYPRJ724EMt5IWmt
kxRM3iR8UpgxaiB+adg5SfkwSPfBNd7z7SRyksVwUwy3yETy/qq2sYzDsIlXMwActtjCs1f10jyN
h/RIbnNJNtIT9SBJL/z9k38d9APUNoqWQDuCVZazr8LMXe/0gb19r889bw6c2yGnL7Bt+o6hCe7c
FgrByIZfjKYoJ2On1lTPYuqYCml4Oc5MGCkmOGRuX8jzbkiZKvcyaofxiG0JnVgKmVUYP9BxR9Hy
7rSNfJFrEB6i3wfEGEvTkFfadeRr3eUjGxbJE8wnLwK7vhfDgAsWcJYyS6ZX1Y1/07jVUDpnAm1v
dKQ8dcGSNGie7SPHdXDNM13ReAnV7J8AdoIefpJwV9xCaMIRmprxXqgUSBKQA2KiwdQsryrojftA
I+Kwu1fC2Kt/VPgur9LwxW+A1FyeL2Z7Wy4OaKByuIMxqpSW21H22wWH5IHJoaNSjDt+/8Cawfhx
qJBM/yUIWii96TwxF1d1TFepX70JutARPeRUbns0OHvtYyUwEh/HA6DSkRyykzoXvR+oJpXnXbdJ
DgnUfjIJ6AK5uCsmfcsB/CgK8XP5ACoRixE5Vh1QKXumwF2VKiDbykUqV2TCYe++BypOjOXATeMS
TQ/6kl5jvZOs/ihd9fLua/eJ1tMgE9JkbgFPCn6/us6SFUq1/Y5eYv7uJERJXlrTst9Um4jS5vmk
R2EhrNKAA81s0amO+6wFG8W9qfS+81V+Fw9KqclUVzmZ476UZMt1psjWQ3vpK5JEuenKD3nohCLo
XuVVrVAt2sC6AavO4We7dywdOto57KliR3+tvRsT+bkpgmbPNMdNt0ar/MespsX74v8cLeD0HG7o
MFQq/J7eTkalHy6c56N/qzMs+isrjbVE8Ad+GFSkU21VITKqjhbPUTSfjidCIHlwTbxvjRoMCYMj
kg4ExggPx2qca+MbCUWLfoBLCBoiCtZzCFZTrokellLp/CMt4zDV6568UTV0aEAtyih45RWnpUgL
UVpdEWA8shArSVJuAmcjTRFJ4qZj67q4USixkvQK0fufjMeZyY4elAVU3rBcYhsOtJeREn9tyoib
26LIN5ikPPt6dsNtnhBsEJ0tMltI6F5oQHuWoU6R7t17OAy1AihSDPvoqL2zwrlonkI94loNFOPV
2a9o4RzK2zjJDx3NllKd3yW9OMcnvklZiXZ3Be5NXnEcLpYaEGKazz0K3106TL3mui8YBXAsFz5r
39LpIRRN7/8/WsNwRcDQwZVDsABFHMM4IZ4D/wLzsacZS2+h2BI/eZhlz+6vDTw/uBQrG8QP7tqf
iyXNQk9rc2yTz+l2hIM/p3Cc6PXE4PTbzIhR2q0XzDEy0CqeKTAcd0yVm59mVhJp/D7tQ6oe0mUZ
U6ioaO1vZwwIGfGBthaMznIzqiRsfEXLDURlWbetlHWj0Ts7YfygOApwS04NMTBIadcw8HoCf+ot
+KZmHY9nVRyGRWjk+Ncu2vvgHn1f4yrHemCpi1MAN+EaSuNgmq1Y9h0pPTO5F7jGWJKYv5kJOy/5
yPysrH2med72ONsbAJbE8tCwNd4PCySGhfnN0QzFEl1eSaYP6sERLZ6nLwa2hk/V2h4GWCZHT5iM
UoT6aiqJNyvReEyZbCaOm0I2vPKlXXL86dWV+Pc+H+5jnFu0+argmlZCDscEbgSiUks6396N2b+q
5xBm8Y3WiGunENhJkZ1cxHtvQpvRL0B7wP+v+voAvyknFADr8pXoWiueNVvA8+KKH+/gNn2cxvaW
KQNOZ8hzq+hwWMLAndC5miKHH4g8cXYuK6zbSzDLTxGyuZVf/yzlanOSPqo70FPI9FyTOgKxrEZN
GW5yT3vbVncVSGS9i1k3TW13hiE1P+93rPU2mYflS+TvBTMyP405unvbKWKp/BUtbtPMBTCflu7l
408sg3W3DmHq8H7zH7gCsXYcKlCqICg/EYKT7G9k1k17FM2+0ZYuajQFo9ZnBZ2CYNYTQECek3UZ
KNpV9EYM4bsQy8wBtDF/Ah9od/t6DI4rNPa2YdtKwXbCUXolFKARkQTRscwFeoYmPFdBp6ISWvHO
yYHNbKaFVCfXTnwEJWAiZ+VRL7qKb+zDMUpBo5P/cwNWfbi+l6A1mrsNsp7QntbMg0eh0C/tKfjV
WLs2E+BJUFIwT4es+12zR48p5x7d1junReCgNk4U3nSHn7xWbwheSbROh1gGWMsswUcH3xnKEMgt
xHdcxM1icrxqMkaMQCkJRQ7kseEaeJwPeo74q6cpDCb1J/zwdzRu/JXzSOGJyrwGdFgf5q+IguIF
aOaBz8+CEqmdzPpf1y/etT6spC6XRnG41B2KUfymDzbUXGK3H9GV4VAmgW782pMv1qId87/jNL0t
OdRtNignl82zwAdVp7NykwlqHe9sWuEf8WKMBVqfuiAgTFPkor5GdzlgAi7gtAC7syPI9FUpu3io
T4eYQ3TF6nAygZh4ze2VSwwXqyl1qtxBpRPUOMt5EcH1dIF38bdGSJmDlQjBUsg4guYfmVrKWp8J
+Zb0cU4ugE0lKSwkWA26NGoH8BbfbEI2wJkkDAE5tEDSNUPmEGam/nhs+cBXO3VzqLPB83ETTlfC
/ldmqRvYNndLVdXSSeQ6VKxzEed4sDTs6ijHUvjDj6/Dg9C9Br/FbxXuxETyU0eg4UfLDB1zY8iR
y3BzM8eG/9K1c0C9EpLbbsX5P/Ou3ntzAYxfI/DI98U2jsmqizhzBbyChzqEyETSo9XQteZh0jRL
Cj8aNsPGYuxtEd4MiN35KUqMSTziMDDg+v05vkZWQWOVD2L3/ROhHPzgYgrfpzoOHn8w9SZZ7yGh
c980n+VIKbR6gw28O4cCNwfY8mZ7vh6gplxub7mNNqzP3pWSXj9dlKY+hH+KTTEdddiPE6+76ttz
yryxsOx4mdSDlBNc8gNXxe+p3jIPfSLRGptRxuz23v7bViGXQ0j/8buVIxOAMsUIQ/zuesd1SRvx
h7asCLXc+DJHC0cJUFkOMy0PlbMcj6CUj2mPIpsNn7g+hIu6n0aAXTi/GVZnnr072by4x79sEP7Y
Na7KoZRdksUJgf7t6gRWitxwpqtqN6yU0ekh7rowglYKTL3b4h6tueZA3G3/ryoGb8ktAaC7ZofG
w4BpPj5jm22oR8HC57AVbm32jGut4PXFNDgXdfwhlPdo4Z/Zj6jqAhxh7GFpyiscJVZpplPzrrcI
TyuqHpQEtbJTWFBFuAd2N6J1/xMB312QDhlrs9MO5lvAJFXWrVZ9o2xuK3SByqM5d9GqPJapdhhd
42uTc+NYy6VCQw85JxTZ9SI5trDWqefsjvI4i/VDueNVXXlLK5rOwGhMSDuwtqFS24dLcVJrHQHJ
C3uFm2kYmYpokxy2Rx4yoJAdAOnsa6RCKTgJFPtphwsQFzenTt0kjkoGsKvmumLmdkpeNGkg8n4a
2DEivJcxvATdNeJprnzuQxuPRVysKnPsZ+Zf1kv4Um8ZE358foG5SpORJwJBPZKeL17shqbj77Bh
AC3TxFZyr9Aqv07wA9iIRtkcNuA6hkGzqK4kP8OYYLqV+RTnaQEkZqlKJqux7SCrtEeGBkKkZ3V9
HevIUmHaAtigcHPmyF3MjqCDdw5PK4qqMrIBt0pQzq7e7U4ow98lz1nh9IwyaFXHMnHQB8gp5a9Y
FQp/c8voPMrUfgiW2ny6Uk1KEP5rCBBxOCZky3aoM02n+e/Qdnu8S1iNYevk0OvHqt5l/DWoIFr4
FZHDenuoH34/wvBkK0foD8DDPo0SViQwHQ4laoUvyaxxnUS0vQ0Ums6egAlQAkTvx0V2Fc8gFBxW
ArMPTiPyBsM3H2mkye0GmS1i1JqbU7hWEyT9yRSHYwl/4oDHnCZjHZaCj0fC66CfAfQohmFF8c+7
6EmSk8NjiBFhYsDZk1khJeWkL7NThzsW1n8m3b37nxVQsMAcE6VJZIQUIHWeSQ4ZEL8joBYBD4bM
VsDxYgO5M16um8tIq4RDz6pEEeJ734CKIyh95mdBqx5OLjGEVApjHOSpSAhMejTucJKwNeMqmO7E
A2s+SE/2zpFd2RLjqdCbZn+2ss/tmZp1ZqQPSHAndmBXRZogYo2oMzRqfHpdkCEfCOQMWcmp0dio
rRJqp0xAWmxzH6J7T93/2xj99Gib++5sej3qlnKhd0Jhl72y7+RG2SwUMx0MxjXoqD1tb09SnDil
egWIIadJOXuxSKVh5ne8XkD6PnDeLXbsapB+l7PRXq8qyj85xKZG5yvMjJqClx2L03HeNlUNen3p
b1VxT/oSEXNF7W/8TzTQyE3mq/kf5Ih/3vYR6pWTtdHksqPNTlRQaygpW7EhyyXqcnqoGkGvDOdL
A6qZ+qcpGiTyTRPuks10WBLKYv2gdSfhAwEPByQhewMHP13bN7vpV3RVjQksxB38nYMI4s7IP0do
vYHIJ6qAWFkCzL9x3y3AsqjYByry/0GV9VoxpF+gb6ZynSZTZGRc/1V1eU3u8eHCeSGQBbT4gFNc
NXgYOeanPxvi26mEVO0REcpuwiSRx9jSeROrlvTD28XVTdOYtxfzHAmwmiUEiz45aQcKUg20N+vu
g2RVVyAby0uDb13qqt4dwGX/bQx6gtG4DIuDppZpHKt0yHds1/X1kW0LYuE/DBihlxp2yu5dgpvF
7yJgV6yCz98AtgFjyFpaEu5vw/whtwhcLf96Iu/gvQARXk619Dewx9t+4ClOHS9EHYMoL0chUk3D
Cx2H92pJaoaIYWgVWSBNKESR5D+6ZPAISZo8j+8E2Y92IWRigSdRjcPFhqHO8TlOvSTSIb62eKHN
PqhiTBgKrr9BFNnNyoy0V1yBVaIEcblXlEagLrX25wuFu0ICxX5UfGOlnZbWn/t3Gel4JGyWamRm
/D/CfINVCJLMv/XguDC0KZ1ntB1NUS1BEUGvCuT+yDNumQU8nEdArzEQ5MBXsQYfxzQxJVfZZFcj
jN8/XPgzazoDYM7xOzyUK+e+Keg737/IJy1QlW0oEXZpadXI6ZufGlf45lGIq760rGPs/Cg7HrD7
+DOeduKVkctuqqr5EecKHaBP/kbgbBlZP6NhjiDQz6Mu6xNZvt93yj6g2KMM+dy16As2mm2hTNfL
vuhSnRxzgljba/J2gc7AA1LfPxvR216F/bxlrH0rxeTL8hxcSrQs1df4+h/qaevTRC/rnl4xwJkM
h0dlexv3DoC99dFrcMqe9sK33y0nxZAXenNdvN0sjZdZiHFP8JgZYVOXX7h2toER0KzA4h1rKKCn
UHJ9q6LUpOzfZSoxlLSiPHLqP/URdEnfBw1dDMtEhe63+1jPqySXrIeI/gDGMCg7kPyqLWmTunk0
JmsUX7E6z/1yvnTyuHuW42iCPqa9QIug1wD9C8I6/wRoZ3Cwa9fvpuHXO2rVNbqpc8FlLNMZTe9Y
5Bw41IfcwGw7ZonmUgsaEjnJRijA9ffu8TZebyN4QWKZegC9dTPYEIQ12Tl8MRnjBoufsCmBD0T+
7X2g9RahxIwaQA9DQRSQFatDFzGHdseQZ0XTdCecRWqoHYgSItH2v8Td7wpkOevXZKr0kNXaUsmj
zwHKDppYmmtUM7MDtjfmg6wx03ud4jtGhGKi/VKl1+7hnKRKAyJaBS9q7JtNAzq3HneelaYle0Dl
QaV28HEv1s7xrz9DB9YtE/LjDIaMqI9EPpLYf5/7NitkfPRuqNzGYRMWfb5/DnKK+X4Ubvtr6Tmh
cpRJZFyMcJoY4uhHRjhqmwYVQ2b/irmzTjj+Edh74TLW59j0/lqignEGV0wjwPIJZTfTep21u4Tw
IGU+cmOkslCbrl38Z6Gn4d0b0N/03qjq5jIz2H9V2znbbOLNu2GN/DcZYR1BOzgQszt8e+qIPwWU
CeAbgJ2XlLuAw3hGrrd+qdPZgt22ZWxhdaHyTqcHoNk8EE5mV7BPjrVADGE2fSAZrrSlBYJig5Sn
xh+E5gZdplIYA1LL2qIcE5vptm/vXgp6DafwqQvvx/9NrZHMwK9yQeAvSA/9XG2iR5B1AHYiu/40
sodcWRwWjVFBjkr9DO11sm0fdOX5eqDAl7C3qgAQRSJamn3uOUpkqzDtHh3jpetkRkRmX8NQ8ZzZ
9OWEEL4GGH5zlyhmbNgwUJLHclORp+b0zkokStrgMLxW9Qu5ArsR0Nr6LlQihKAc3FBpt8JTF181
oERJBZyS5BkVCLmT/WzwrOqDRXZMDzaTKQ9gUGkqIGJi/A0aCdZmoEKYZ0Ed6YM654YRhghZis6V
cfUtFek24vH+PM9VSeeRgaeRC4/vDs5Z2m0mI6aTSCAj7/PlDHcMXPSEKFySTyVVsxQMx3772K3A
M9qck2Kq53Ok3fHZ0WSn+C0dKgvVBxyXx9gjOFGu92RritRYb7rpfskpz0zruD8uBvmcjC39wzdE
xOla/q+XJ8L+h92TOgIzBzkkJAbgMDQmOm+rpB/794+bCIGCPYxGpSdPAgSJMcBQUSLegU7Ly/B+
WNpwYgfZJB2OSJ7mXk6nVKFJgfh4hqTOiF1Hx4bCrRaM+p1lR7Wvcu23pBSlejy3UbTiaOVC/OwG
zC3OtU0eEaRZEpd0gcocqX1p3pVFU7mm0Ub9NjZ84g7FLgX15YnY4mwgZkcNNxuNYOCdKtUIHFw7
OZo81oMrL3WSUPPyJgyJNRJ3SqDTs5GjKKdvnzW+pZGMRjqGQrmQYI1pS0IlBu7k1LMjxgy6TJ4j
udYaEqMCeSrL3Y5cI46AQdFKTyomwztssLTtx4ADMXQoDItKZdvvkb6b2MiqhdoVzveeaSJLJvkd
vjkidVYOcN9lWA6vYRvCdk6ZI6CzxfV5NvsoZHkO3kpLS7eyi6pHguvWaoQiW8QcFmfkUC6Epvwr
Y+BACdr1QYDmcIkJaIL3ThYdxA2y19jJlWvTeF6NaJZ1fk8Zzi8KAyuuCafzJ7zLYhVaUbgCrTkB
WrD9fc0NJDKWwCOwOJoaPP5q/AvDQma/9KCLtkyTHlj+mb//GRI7H3dW6baK5Hysd/kJMWFV4fAu
aXCHGKZDrOe+hlIu/Bz1DXccLWaAMl+1eJDehWjRxc1LHwKa3BQOLnXJs3YGzrwemqJG4tfRYqd7
ND/INcr9c4gta7V4rhlkAc1rzCkguVOYk8CcjQh46YPXfk+bz6g3cBIwbRXppZmWI3hivwW1LgDg
/53moN+j5pTrNuEOO7NUp/yGRRkhOkHWq4hgfWilfBp4BpvscprdtHjjqZMlbILuWomTGMxi3p1u
HmAPDpdeumOsESaEmwJQQHvcjBQFVM9dm7lpwjaRuwhpl5aemhJjYfNbSmieIVB7DYYK4x38BGAf
5XFAxyiUtHq8QxVsjoeNWB+r5gPYCqAkW167lX8zedVevhmafRWlnZKnQmLChoQ54xDxtPxcneiN
YX8JzloCtRXilWMFAn4SfZdn140Ai5+QVG3Kb2J82ffl7jsk2/urdz+HMQ8Tjakbo2hyOvqOtGXX
wmBsgw654t1YjOs5Qs4bJpwBfbu2PfaA64esyFvuOWkhjXmYgnr7X++Je6ODRAm/Wmnh5LNZbiOr
0DTbHykGxsSwSQvKWJILlWkHw+ARwEEzCAVez5evgtrJb3mResqIxGqtNzi7VLhu221n2nJS2kfX
LPjpjBTpff4oRkHvIC/f0iRdJVDjJzq613yTkj32t3PnioWhCL88GcNfdWl47p1HDx0YEJ9gt5bF
NQiJrA7oWeUyRAaMxmi3nDv0HXcMHQl+kiUAvNId14hWWr0lsOsDlTpz6Swczkpknu7kkSTdYOIG
kGqLH1glSROVXjsTfRgUlchU939759BcFgSlMJot+U7WImtZ5EgO2uUvezrm+SIpUwmyfyiCSan4
SDfUH25d3uUAFpMZ3zwZdthQT09gBJdEzsFZDZL1uF3jFCW0ehcWk4A5WlSTrS6Huzk/mEv0DQqV
/QF3r+2y8z2AcGQJZtTVRUOYE4z3hCLoS7KTLUp6ZkrPIea8KpdsL3iLnAeCtWfukNNkuOfir4F3
MRa6HJ/91H/Bqr56Vaa0MCVn0vGuZ3fZZZHAqKZuh77BUDu7FJlNo53w+TFHR1hPVwUDoA+tK9IA
W54cAXtRtg9WqAWv4zspuTBBlPiiSTvltck0ng5hRGYLt+1UUYHuubhfX80U6h3LyPCVkNVLft1h
+B5hbt/Dgq4skNrJyweY+tsTVK85H1m71cixHelEhc6fY3KLSNYMdUyWD8p5dAmlMDpbz1A4TZRB
Xd9/lr1wlLej6futNDQ1ks02YFdgP0ln1wW8ISDEhQILwg3dAoojQk7N8fi45Q0QH7dDx/IIvbeS
dBeQ+KmDbG1x6ZpI9zKHdvH/vZV1UKA5/T/9I/HKNxDuFOu/1oyU5Io/GDpeqOfDjhECJJMqw9Rg
TAQTyMr4LNs7T+48YxjXN6V9mDEnYElB0nK9cjs0jo3nD8hyfFB8zBKKKMKbcvK/d+kaKZAQwDMS
Rt0bVnZB+bFFpYrn6V1nZ+anwlvYNJGWk49k5ts6S2iPU9radxLzMTWCY7ba2LmGVK92zC6A/N4+
d4Ur1SRfi/n4W4FLdIwP0S7a69ZMAL2yXn9tKWUB3Vht5xfXbm59/B2mev4xqqHBU0IIFEawdold
KCTAPc1AfdQNGpAKAOfX6dMMjdHnkcFORdgRwuD86sQE9M0DjvRRR7xnmWlRUg0LcUNmqGRPlkvv
aC07/BFF2sZqzaD5npbqc6JC9UHquqc2Bvw9oXDCgKcMDPYDNGYYD5N5e3ZUSaVkf4A290ThYBnr
+bVvSVU3DRXGnSsCC7BndV8UIMsLG8Z6CtaSMdEl8uZgRAhDS1+8SDScVsW/wPVHU83nFeehzL4A
JpKpeCqWt/JCeSc7nMr7ya17D7ss/WiBh++5De3oXdMuESGbov1QEobugNirZQTl2BfoapLOdtwA
cp/G9xpgSmTYCEZFhOoatiWdNpu4NeDw7MaHnygbgAlxk9P6c21I9eO1IEpQl1qv2JjZLNV5+z3V
Hqq6Xuq1YhORg/M8gisrAZ58vhOrw0i63szfqUuXrRwWK9vv0jUG9NVMj2655kYbvW6lg1SLWrHC
GqbpxUKF639zaiVUyoA2jZlF491Co48l2mJcmkJPqVSDlck8fKZOOCjdDPvDgZU2MQ7bTkKmMX0C
SZJCQYWmklY52KPdksuOYI4GSBvIvOx8dWN6TVYcbe1+GEbvn/8YiHGhb/TkrPFDBwVo24pCvbsz
W8f8+r+KOcKxwpbXQNgsVeT+C0f3QgOQhcFgUP1ownxeOmPt2cUMWMrYuY2vT5Gm3XDlx9l7Yj/v
vB05rNOGcgipHG7l7d3DzjVP4y4qMNJ6pd0kKfhsHHixtZRxJnf3z3aGGKLf8RT1N4FTb4oiD0EJ
BFMEWGgwoTmK8HIpdy6lm7JzvRqjEB3S8S9lAJSrUjtvlJNGXy6dbGwqRhaBB3ITkj+x4/rQr/mn
PNyFNm4JAvvQVv9Ly7fTWxmh4YcreltUHxZMAOWDtU/H8QLmERPrHmZnT/n3vHCNwyeb3zw7Cy7F
NEjfW0gOogDG6yJ4GMUTQT4onnadVQXrJ45sYxgGl/N+I7VXv8JOuG4kCXAf8XLXJLE2vxbVlqNE
3plPKHk8rMiy7RlT2I1cNMLYP2sTpyNHjqjffSBQnmSbcazSntd5Ylws42sL8jwDkB9sZiQZlgvv
qep+NqQuSTlP/ero+7SFLF4s4Eul83z7kHSOynKLRrZTDsjvH/Nrykk7t1sTxfOBqYOryXkc6XQ/
QGlELepOP+P9F2NDC3QaA5nBzXAJyFH8Y9QanCMyRgEdDAF6j+XFJW26Cv8Xxcv6dlszaT3BnBlZ
s93wlqstef3iQI8aAZ1b1vxlyf8mG8M62SzYYA12ur7r7E1CFFD5yAbGJa8SN3fQqUcyiwPh5IUl
BXG+pH7Xlp28EamN9Znx6umRchFMQ1DFatCJoIDWo8vN+I3AbRW6MA17evGGAmdusda4LtLQcpFc
l/0+kmjUIi9FyQxstpYwvQxdXbA026lyco2FnDRi6XYjULm8OE9Vm29QCsDsexgduqpErcsPDXRI
i/l2s1zR4gNny3TdEpMrnqDAxDSeeGZ5uM83avE9uomjfk60rKBrtkAdQr+Vn3e8tDHTSWFk1fgo
w6zhL0B4abiemsiSSRCWUu4a3DOBDfFmw5GIgQ/aWQ7Vec66kEUrbtn6vPb9vFP1rIWZMJM6uYuF
kZHgubi54k1HheA1dBGMCZXn3MZ8wqBMdoO9ny8DQhFUb5Fb2whb+LVBCuM/xUO2fWwzfX2VQQ/A
Fg8WIts1dhRkoHeefLlTRhqsClbN8kNVe0puMl1BYWTUP3UHy+/O+HRJy3e+bUiJHFiUJ2Ikwzee
OZG9YiD6zoKvUUJ1FlbSFnhXbD0O6DnE2hc5DaoI4uzUm7q+oMmImLOQb5oT4SxycLETHzMcQz8g
D6Jxv+BgwLdUPHvzmD1UKgbUSzAsju5JJRSssStDRLf5+z/xmlCUa5y4YkIeYOmWmyJqNa/ft2N/
aFi5wlYPanPEVhdRIm68aOSg6ybjqFmVqfs2bOazPeyF7+DB8FREFEzMNNikLOdsixXqp8Du5yae
k6doiAxXimINAqrDoLBwIK6JGr2kvaOAUrdA1qwQ9jvSmykq8u1MuygQtr25Ng2WVudL7NwR28tr
yn3iFMhbPqcRiIX2HYcm0YZcP89UC3mAZPm/ICZd3WTwYDBzH2j2UDerZyDitPOpUYMZKY1yhUBt
3eo/Hr+KUeG8g9TP0ELMk32p4P91yzh4pIYcxdSgKpEP/g/MRDNk6I+z9tgvUFiM6EBD/Aj21cun
t+qIfPsClnJ4NvLrphdynUWo03bsVzJcPsev5A6ze3L3v356740Tn23+054na4TBrBd1yDTbcau5
XpqQVFiPoHCDfPA2ykj3yAfBZ7sOboLxAi9dcPqx/iMBNv4ku7BykVjiVHkycycKgWwEFIYefxa1
91Kl5xqxomo8XI/qTSNCGeXWKGUG/yCdx6k96ciMYq63iZlx9z6KgPP5OAbRzbiLU5jZJXmvyL6g
qqd2fcoJvy+kPIq7cB7Eg5acrQfD0K7K1uXkWOPIbPoLsbd4BFgvmcIWPS8/HtFA04OjnuLFYb4Q
Ucr84gkIvTJkAgmH4BXFm7vQCyBCYPS988bPrDZLkUdhSFfWB9T1xaZ0bq9VvDvKyryaFtBYF9Su
+myf90B7w18Nl7OuUXfQLCTn3KFG4nuoZjYvPSscdnJobggxaZnJD7yAmwSR+jUVeYuJg12+F9Rb
piAELp3n3urUUMPRkH8smrUTn5Bwl087XY6Eqz1o04pm6fav7nE6IRAXVkUpZ/V5IG2+TrrDgMLG
L1tR6MazUbNQJ3u2zhMCCklv/YylOd+v5VwvvqrQU1iar71Al3buuoBVZBGEtfPalPpjznjEpjKO
LKtmB+kThn5XyYJSULjfndO79slU88eJysmkSGoPxHK4EBBn3CL0gym7tDKIJAVjQyTGNN5mcFf1
1X2zxLgmEloDFkOpZc4n+GL+mSLwslEUo1aquhScCgAPHSgwlL1SyattMa+Ul45UVr9bbzKhHXXD
vaMNWCNby+STVlIZvBUI3kJHpsjgGQGAClwHPP9qwqGkbZ0OlgYgVudqdfmCuL+USZd6dU+OB1n2
ygJcWaA0t1O8tPhnJoLyN8dMNzY3vwCGsXA9yzJIb35Yo4coPo1Q8Oa8ziRnyzPeFmmGt6dpaJal
GXXuRnuM278KCG9zNdZCXGLuoiubKkDdJOM2o4id5Il8Q6s4kycibzazDSVZRaaFmLDQh2EiD/7O
+ap9Jj3vRjXAGBpHvnod+StdpVJV3wHFvkPWT85TJWmjaR39nThtnXvMSm9edfCVgk84Wr3493IR
SvEEhOkdyDSDQZI70AFbwO1O5OexSpuER5rXvzG1JSp9AuWIuJAea/HkSd5ls2A2fXmoQ64+WOvu
7cLepkLKt5OlLtstg5daGiepQ2Wx9cQEZ6mAL6eoZbEXgXGGyMS+uH+7SOPbocaF1Szm8h5ziNmo
5bZd4u6H9TtJ0rESiQOUZ2LECYoLFlrq8fTmw89oxM3J/c0Ppw2Mqbz47W2DPtzERBT6E3CZNNqQ
d1ENTYkScKu1ZEypo8Us8XrR4C2wouS4p+YrPYPa6vl3yq7DUeslM1hFivJcI14rkcMDg6ej5iC/
u/yVAgvSB8rc4/66CXUfmhAS2eGDE986SVb8FfrwCl4w7OS4K0xVVWN1NfrSkSc5PUSxANXaIPhS
zdDlpPgSBJvNf1H9YzUCARsZXNPQwXKdox0VBNK474V61rvpc8fZhuVYnxrd7vpGQ/3vus7D8vtG
92exu+cmzF15wnW96/LQwIwhWQKASNM9BiqLAxMWhuB4UYYckRMibvOx75esvJS1boWgJmwUPxxt
biqVp93cmqCyFXxvekNrQEhitzL8czQihhfpL1BLPlEiaWaBKztpgCiXwNzE7eBUcBGoXis3mXhD
eZ2KL+qSMBl64ZIjLhRzRD+enELOI9XxvMMrC4bLFywzXYy1QIf1Nsb4CLgo4k2Y7pOaJQ5t5DZw
5kEXhcXVcS7qBF/VhbocUmlES09K14gIRoYWBLZGSF314KpUh9dwfpg/yqH4WMbq3piTgvNqAnA7
PljCg1QbPmYpADPDn+fc9dawJQ8wCC44L/60YLwf6oNVfM8n0kunl8Zdv/C4E79f/B/PdLWfJDky
t+fmIy7GmSnxnBA+huOtX2/fm2ZRAbOlHjQUU2+xQCcT2PO0KXiFILXdE6ttItlKSiZ7q2C68e5L
f48H6wfCeqq69uwP+qHeX0v4/7uZNR5S49tCivAimpV3GehU13V05ctDfaIX87aBmJj7+5Sil7Ga
1NvkbqT1femib0kQUsNqD5B0haP9WcqB78/R5VESuRziUk6P3qPvS44q0i348sU4AgY22lLuoDf+
WJ267MOcDBaQaqDnM7NCSa5eOwyMiRLIobpY0JJbOmriur5Dttpu8qbQq8vwQilN2GdONMndzyzx
OI6lqvLaE1oHxEOU0G68q+ld7b2uv42RUkD7y0w76BXzbA3/EULOsRO1MCH+vijREac340CHfRr7
wS65o2+tG1HeRd3InmPVLwtowLvlkFxQLRJPldKFDFpkwY5H0spZEPb2mM+B4k+2jfTgy5SA/y+8
FN0NzK+v+K013nnF7Vhj+CMKBdXjeC3E21v7THMeJrl0RREadW9Gg8J/ORyR5gHOWhHXIoLJG7us
kbzg8u1j9s4B1iZx+nuOU7WHQ4jTbkaokq1a/ajZJsQR4XRJfex7PPCR+4hHrIMtZnw3uJERNK6q
sMvbWTBvZdI+GQbu+9umS84EgMNJJJcibHwfRL0B/MWN05tOsi1io1aivK9JGxaSRkNAtybG0Rk/
5xwfRhbK/oGIoUdERX9+Gb00v5P1rWSivnZCOpxSqj0JwT1OCaSek52BrG3eC8D3RMukttn7WFVA
mVDE5EZwSEGgd6R5CnF57RILJhxIFtUl+6cgwWG8qmXbAz/TccyRnKsXGcSlNEgcuvIZ3aiIuReT
PNVagJwWwcxU1A+RLB1HA50qy4SQw2463nBKwZ8ixP196n1Ga5L9RuRDC5nnZ+375/E2N6RD6uJr
tY6YTolUCum3rLuzGspTJenR0dw4gAlFWQHvzK6xOhEXWtRpqbYs3HGvWqUnOZirtM0uqHAUnpoy
b4ZWwYPx6NMMo3snWPp0cof8VAGWebRFsMDT4dtNfrFxO38VLmdd3uDb6Mxczicr/3ZabIJZJgAH
D0N4A3ENv1ioWfxFi3Nv088dCwprPS+02cy7fALZXWAuMZDk7vehnFOkFbWxqHHoIjYmFhm9HTvJ
AAt82xuo8rOZtqVH8PuPTtZJXyQIIt8DPGmP9gyRnHWxDtgplsINtJA0aNzOUmkhcJJbKNfxOAWs
uh0XK+WWRw5AzX6ATVCluwXACuyMZTkPK0qlMo7+9aNtYMz0zS3ASP/3q+Uw+5CmV0BWzw8Sjt/T
pQDN+cqxO9dG9YY5LmCH0xe1CwK9kQIVDcr2J+TTgUZK11SiLamQAygek8q/tSGj9TtI+JdKnNIg
JRQkQxDHcRmCl/ZpqBWSW14h+QIlYz3d5mlsS8Xelr7dXo+msu+sU0pxvsImDj94SHimAlt0ItNI
uv0NqVeDnY1s30WrN7JBESOSk+tVBLyBb8xwWrREELV/tbguw6b9gRM/axxvJHF8GSGQFhGbc0H9
K4Ee1Y6bpabZHvPKDn4ibsYSjTIondiuVb/AYrXyGo4G7gWFyQl17q532/DtwVNjFt570rKIGpqf
3IFTlrRaU9mW3oOP6JwGeB/2Hz+Ya7rmjdvlm+eApPYK5HSKvUxLQtkLUMaaIrVT3urkN1ecxrZt
POrh+tS6hzxfqU+tmxdQMo3TFCJGPcC2/95tJIDG0fO5ybigAblvN+Vus/1+S8Pn51itQnFd/1w0
UI2rnAMwWqJVrdVDCTz8IQvxT1TBMyBPP6IBa6uK+Of3BlvClUs7BnyDDtkB1IjoTkb8I8NwniWh
qVOx07HaBGRexQMQ7QrIF1PeJWEby7ySNdhEWAFWopE14rvInuqsybPt0F3wJuLlNNZBDXFZtmqe
UOWWoPg4GVIK9BFHrUwhUgp9MPqWIpwVMtsnkKqugFmGkQP3cDBA7n3K4i5l/zoxtKm6s20f/JA6
/INv/wcGm7vrae/kC5UQwUawm1VAYkUS8wiSs8y24e0uK7Blc4nqi+hnG3rIa3Wwany7W8SN2Fkq
BP9SQfpyQXMdrdqRWz9bVQ6fpQmqVmMNwlY1i9E8wYq/ntj3BS2tIwC9JFCvkIzXrOSk1tsxkTNt
6VolAFWVzorVOelRTQ/aNAc68WKXfrkcFWdcJ18Y9Xntr1KYp7pH8VQqNMSmoqm1aZ9uRxEARPy4
TUFpDs41eoIWT5osnSVFaO/YKhwgs5f4013y2JEBYsl6wFrrl4DXO/AmE33/2vZ7ZFdc8P9cDiu7
We/pyL5ze7rHFhPVKZ1m7ZLkuAvfbQRYbvW2vNdoybfz5ZRWZKjxP3ZVQiARJ4iAwNymO2FklJO4
oFh30Br1l7iSILyJoNkkNyklhVpP636v/qIU97tlpFLhKKVz0GqFpBKjDkq/5uz7fyCq58kxGFGg
cq3KgyprzprJ/R1Um+gKy/0YxZi6maI8e9pQJ3mBO25gW7h9jg4mTjr4h6g+mNUbcMzqMrWAPmx2
pf3xSMIn7tKU6V6fV5fkX26kfenKCt1f2dPb6kh+OmFtsa7hKRvSFExuU3x0KIQdh/sX5fpCbWrD
PuxOow3krpAPQ04hI6BKjJl/XLD+GhfvPs3MTCofy1f5IXEtc/1WeuKALALITmRBC0n9daf7Hs3n
uWfWDdz4/FfHc0LO1cWRR9bwKJSMGHMFfHSp+basOE1YJ9YVO5q6sKkcD3p9lv0PQ911gR/U3hTC
qF90q5jYPLzBmXBDTo3kvV8T1qbI2aZrSkbH7qKyGaR+oJs29wvXz3RuevemH1bABMHk3mSlY3DM
eNmqejw9UGjtdhnigrcbzKXOYG4Tfr+TDoTvMvrr9uvPsm+/GUXinGtOHRQD6irJ/nfdKecpoQ1Z
4TZ8Le8Z1NruStFxdceqMfQBzgAw658KYtYEG8E2UYvOeQS7nMr9lHA6U5Lyku8CmlvOsvF5D4ac
5nL1N+RVhHLb7caipc7BPFsAEqyPC312czUhmnaD1klCpb0IdC35JdnzCRG7XQAE7MexZJCmGucm
K9mEIjWGCHZ/fsLUGECGZ62awnUYn2Q9gafNBgOmUv7cqAhtaefZrDEtneMz642Wxy9b3GNg+J2Y
gDVuAEC3TT/UG/4y8U2fCYKwIpbfSKcIBoDFOvXVhP1R1YvwMMBnSVwFZTilPWF/0BkAWiIiJ1dz
c46z2KdACzSCFz5Cbpyusc2NMx3DC4j8TYbEiesKaOaggObVcipcGq8UPihJwbQeNLXSI3/UHTpm
zfK0FF2jz8A6If8RsZu2WP1uVq+3JQr7UnzCKcYpEEMrmtwMn2PHzjFARNF26Ts8WRKTaZpw8d7m
zS3v7OBzavOlv0U1KhJdLCLvD65ryqGAEzMGkrjMoTvYLceEDVmhK41KGbj3xC1PZ2sHk0wUQI/c
u8iKZOok5Ni2cRSpDOEC3oj+3rOE7w48xNfVG/AVL7RRnYzLtPakWrirgRrmf35IPhVGbP40/jhW
QtOT3QggBvO+T70vz7MPKYHzUbRdk772waufXDTlCarn9Q4Kw3mUzRzL65KwRW/jhMxNhmTcBeIO
ZS9HNIzw2EbAbbUChJkNU1PL9kwM4aMemsZO47Djuh23TbjCvIOiAzfmqBuwhO9hASgn7RheHrMc
8WWyEPo83yihxxyrxh162jyuf68LWZqToy5XeEmFh1lwJl3jXixFS4eqnlseHxz7bqknppCnes4n
5+tCGke7wUXNy+Pclcrd7fANxLymaAff73o1T6r/e2LI6jISxpqtcWKLmeDbPbH/nKFcnJtMNPxN
uG5vuZjz17UZCh6y1Cpxs6twIYl1afoCOnpsAUr2dS5LAn6+fD6fNNbfn408NLDMgH8KOJj5OQB5
MUXO37aky55nfG0f/6Zc+0deuQYOE8+Ci5rJ81yYusUoho8azKj+LWT7YFn6rJ8w9v2lFvS+wbiT
0T/lpDabmo4v2OSLfC9bUk/2vyQO970UNG+6fDKk4KHXgOlCwTIzP1lHdp9Y78JW2RJWEY3MaRie
QvCwBEG7BY8krgE2qU8/9NBr7Mz9ixgtBL3XBsowluoze+dwr78GopexGfBmXxQtRqxNl6MYKix3
LOxAX/7BAiQTLEt+pPj+E6oKMF7fukw+ijAFrSh4NN1Je5PWlHCHLmAnc6DU3TRB8cPd+46hUilU
KlhTbUKIXOO8nN7IfWeIICyrho/UGLefNRHeuysLkW9FpL1aYiSv4QsO2lNOV8/KFoh8aj2CM7Oe
NFgTogXIoYIyZEfWV9mTtVbiXYNhfg7Ef+UzYsXzoafU6uAiXFF85LeDNDeyvYOquQIZhHW6xI5n
Bs67+aLBB95QVPdIzNazukCOSLd+r9uP41CCjWP5WobDwLEZiupVFM9FqW9H8tFWwWKb2WqtCBR/
Fj+VAzS5LqzDGQuNyJR7/I3Ujs3u7/ZSeorw0zehepHMFTx07e2YjhwDFeace1LwaQGaEC6mL7HP
vdGykkVCuwIByKPlRvjoH3EvsXyMCCKGa3Wq9znW2sK2RqYPOrJfE97NYbiS4TtuIYTgFnIx9VqN
Bv7/FieN5+cx1RGuB1cv1vWXq5WRmt2rKQJuRIManhMqjy6e4nRerB5Gz2zMZDOMtXzXOWmv6tcU
dB3fkTnXospqs4vLmTTF6TYrGGnHliQstwADZpklVyaDFvK6B5Ik3B6a9i7Mh0V3h3PJpXzYu2PP
7EmckukyGwExAWTMUXb9wPh+d2V9ONpR0WE3rEuq0pxXLO2K43je+xim3ln7jm9YCqNzuglFunQA
InYFoKfLMc4XfrtX0witMfvPLpyc7+41hASE8FZbXrXPYb78Haat1yC3MtSsk76q0jCGVHq2G5v3
QZQ0SFLch1sPdybTtDd9moi4aI7Fr49yk4g8ScEohEoGqpwQ41QiQcop5g+JPyGW4AsQ6kvyZl3S
qyrgPHKfSXZ0MAV5Ft2QilvHBMGE+eX9nbZz1VaN9LBam/eDn0Wd+2urd0bXqEcO6pAx7Gc/4/MP
5gIZ+w96vwZzAXBaB+Nf+8pNnycyuBHdONlZweBNQVgdSb+3KVpHp6TJ12+B70RtXIYg9x3t1A+w
J+i2Oq7LRA+jybzuJGrYlJK/3SJx7YDMsUI3LYOr7uuTqAgq4b7PNndRM/r3v9YnPsneP4ctndvD
FV1UWv89rUC3Y1CdrmH830xF2It/55sigx/4ui4L/Q0dmfYUsZ5aS5L8Pf9uY/94Lab97z605K7z
6DRc8Hv3KIZ8Oj5+hat9sHIc52Jd6i6mhhk3Kpzd1LkOfUjXtkknr/X5ySoZgATMHt3QujzHYwjL
UK9dNgcJ+PgUQ0mOpEy7mBBjmc2PH+/71QBYjNer9oRmucBl0892co1de1ZzcSbqIsx5hc6xCm3m
cCIuYtJ4Q6vpCQjhB+6sfPgGPqk6UaD8JcnjOmO+EldffgyTmZWE6S6/EQhKHBwu93IJfm2KnNRM
K0FV0eOD/fd9JrK/waDwHXGmZVs/IFqmzxKd8rgbAscdYcZS3IhmevNeUvA2bTP3igBg/VsJ9K1j
hh/vDbPE4YRziu5c2+LjPysMZO02CIEvCU6CAqFbmSbykAGJqtek1SxTjnIaB0Xbg3XW40Hkpnv/
iD2uwlprym1FoshzqmkOdKwnDIyJTew+WOh82+BEhWy583Os3jRsAPcxk3C5C8/mLxeptJ5ZKCs3
S/2n4A6ANjptehurnjf8PHKOvAFC5bBdk1v81YZl2eBrer68JTIgPmnrKYOhBFMVU4ozAVdjA1ty
GeyqXnLtk0luVTyV5JyUTavJ8SgJHzb3hNJTZYd7uHacfCR9vWrYjelJyV3tdo1mTR3atlq77hBB
ykW4WRUVYmahTGwkCvMifwCxBkduAEs6TwGHobNQtnoG/7t2MAwxrHF/gz2FLj3+p+jveUXAIVwt
ADy7M3/cTGwLc+6hat1Tt/kq1wKkOW0RTK3j4r3v/TPZB6UPME7heOifYngD7KOwVKjkPJUfu3R6
u6BMROxHsdZV/6CevyRnHIecInTtD9x0T+Kd2lH8egul6+g37lS+psDHKOmiBfwhqbH+Q3zKyjp6
6nn0cMXQ8PYxcH6ITqO+JCamjd8iT0iQ76lh8DMmmNhqlXN8VmuqHA4MfSym4qzJD3w6QWiUM0+s
s5AVKtLrZXcihA9Jc7z6xObSkh1QibNTRN81AsBc0mFGemwS5CBiGsRXxGI1VrZtvGFhTRz5HGrH
C7UdDq8jFeyAjcaJZMJnaAjutBztRjJHB8/qOJlTI+8W5gq2ESD0oFiHJU+kAiH6j/Mq7dFy7Jx5
6Q9OMKKA1+CEamHp225oT+4ynr+blf81/nv+RDS0XJcLLHh1C+ECprznO20GBlfs4MrTRp5NvU4g
AeZfAHBfvEYKvTVUuRII3jNPEw1yd9EwMnlLUFhwLTWUcgh2p1EdV+NS1KcHOhxUZ6RAtUMpLbm8
RiLkPIsC22VKB0FqXIcpsXPfjl0H20F7+1K5PImTbW4GudC/LNrq+hrutyN6ilHtcPL1e0R4iCo0
EyHCrGzK6RA1/ERqw/fbargG/saa8AY6lLhBDL6If8PyGlK2w4gtUeUJlSTISE0kkOyqgTM/hzcA
svYZdIJDstvmA+vWWtIz21f0+Bq3ogaqft+5SYjUoK4NquNFakYdm7BmUfgCuZPwbYbbsJw0w0bz
47CqkQgoM90m8E5ZY+oZmwydDzYw2LOepGSZZaUgvYZ5wohlrTP8onX4h8pwlfCOu3zfA+43st6I
2kldwHpW8i8O9TU3seRnQH02zqvbCcbdP6hPOE12oAkVlSuwFtDt0/Xes3RpSaaj43JDdVC3r1TZ
2y3+zdzdAdhVK1MfudZoY8KGZYYIoUQ9aKu7E+ElveJp1Rbozxe9ot1vaKx4UVKSOjCUjbxaYjna
YoJtsMDaA+YZ8Keh9VjR44iEnWn5p/HD9kO5AyazHP0/63qgcb9XQofyvNqw9JEgRHVzWd/34L//
tuhIBg9TkOUyDuHjRf7ThpfExhrx8kPtPeniK4rdENFaeGtBDDiemIabksuyn2ihZ1HoTdiXjV00
jvKh+4XRQybyazrgZM0g8DaBRTVkmAVT/hKta3YcBcC2VMz74/LqVjjlp71XfeTqpJ5qrA/u2Zf6
trlIyS8TFMFjk3O3eDljRIO9m0p2Fu4Lno7oRFYOsWt+RsTtTDz1r4QYvmjwCVyXhT0zVBrCcNoX
WY5aUtr8LSL9CZ8AUSERrrl1YE7vvtaUGsJto4gOCjdSDniO/QcejXYnfl/RyTpo51yPPD5o9qbo
kP3330QHc2BxzROGNXgtNKZSbD1QTGQvgxp017h8MhEFjqB7+mRESU++cfY91ntgWR7/JHRPfBfK
ijZKD3zOjGZ50kha4Sd6RfQ37O+RDNI31VmVdh/ulCjSQjdgwFUJQJwEDKyh2uM/W18VYLFaH/uz
h85fK1qozGSHlwaHumGJxA+fFu88liRLR0U/VVHtLOwMXOch0B2fbv1kMWIQDfCNI+Of1SrJqdF4
Hpss11YkgXxCHq9nmHvrPs8AsoKTdy3nMAUTgE/QSY7o5v6/55tJfCs/ncY09k8o51o25UUlaQRs
6o4eS29/qc9IXwt4dotfpbJ76uAlSF5eqnyDm7B5LcmbsozcAiKnSAJtc2m/0qm5irIQ45ACVMC8
jJlnO34saxXoiNUJYIJ1nLU7H/82vqPxi1+NeRaCHJuzQIxSx4jO/AZVO5YDfG8gzaYgL28Rib+r
xR1z8Bm9+P7T3K01R8tLabALzCus2M03UZf0/YlgrQLegBvbC8pQqwKx0+6BrJwEJkfD8923q50C
FcP0eZg+8UO4EN28FK/pCfowz/bDYl6uMBT5Kq82LH3imZAi76WISbAMxsJ6A8YmKta6kz/s9rz/
N7Ud+2PwmXf2qEnOkfSe5tBQtAtV8KiABvLe3Ahfnb9K+H6u5zMXfkWNJUveNnF3SxLLrE6JM5BA
JvroplZRdCIKcYuMjnAz3ELL0m4JrFt0/5hCV7tJcoVHeigoEdQHADlKO6LiWlSwmJJ2iztk84bm
dOy1XgujGKUzL91/mesTUBT8gp3usqXhthdTYjczd985lqa02Mt4DK8I4SfNmTZ+PSNuj3kdfJHE
W8kCIA/KccA2te/q6P5/hsUtN70CUqYw9iV9ZMiFz5JFF4tXKzl1Dp903uYmLGzLoXOmMKxP8MmJ
wc4JbqCiPbs+taU2k0BC2XOXM2UwCEd8OoEcoO8ouMg8ywa+EnaaKxsdC0gdQG3IOD2O+fig+sgB
tVABbQM2ptmFxc2ACoGlRNRT3UZX8CRZk2P2M9nB1csBzM8Y4G1EqQpwZuTj7FLExzKCxAHsckYR
HYSPrWa4rotMLnSqWcLAcj8wMdTCe+TIiI0/ocLIyswM96t7JUSyaPJipay/asXxBPz8NOrrS4mv
5L7ScTDA7BF9EyQHP1NC4dFTWOTdrKqzQ9HKjO1s15ZneC+HDlYqjqKfXzkAZKnr093zJKJSn+1T
a9R4O3e0CqXrjS1ZU51VmwTftgdx6lBqsW7YtrJ62uO15GrPD6nImrRqm/qhtdiUTvm/8LNPhMmq
F7diATPEVUYj6AxEBMi217cAZVJ/Q64xC13D78kXgrbJshcvHLItO2vD0cH7lQzU+9o9OwokjtGm
U0EaVoH4HadTI2wii1uykpljFb38ekE8ean3cewwDLBDgGCW33N/XKYuz23YPt473EHf/1MVSo5P
AGvYNYE2O7SoZVYz46w60OJrVcFF9OHtsPmuh6+RSjIEaTqEPH2WrRg2AsHb2CEQnRDOeTESVFHE
7epDyNW06b5ZsHafpmqG00EiTPJM3UF8AzYiCciVPs2ghPNY/Qwx3jVRjCFUUBxH8ctMjA4n7IHt
aJ8zxO+4cn7RbaQYyGI6C9Z5fqvwnkP6IRI4/WS+LJLwloIWwML/HaWgxIb7q344I3xTYiMRcX7g
oYdkmTGQvWeHMDzlEew9gS+DHwLOdE2gendM9u8J2xS1H/OeeTM1HIXEvYcHWrL0iGP6QnGJoYsL
VtqbDb3kZghxo0OBqOfVnfesxnp1kntRfyW39HEUmi/SG2CSH4VHUb3S0YW5wep6wmeOqWW/5u2Z
5TU39pfOD+U97okZMAc92JAi6yF4k6CSGxGr5RmEPdcYjV2ryjrkrAltU0aqcaXfe6e0zcZ9N+sF
JcCVVK/LPWF5H/g5H+mRGs/yAPtZidnqEfQtr7VKRJRIrhANIlv8HiqvJoRl3AKJtbDCML+2V9BU
9P//jLDRWkwN7HesYdvv8x9R0x/HvJDsrQ86WSoVzt0ZcW9Vt4q1jcYDYzZ0zv3DsjSb2Gi7qiDp
HdBC0OeIqsAPernqg9XKnhxZmwMDiwkFXsq9gtY+nx7su9z46WvyNUCMnrsjDXveAPpdFEJoIAyj
Jbk94bIhINuRLBG1PFw3hNeVFaujtDUfZdHHKdAojjHX0qOaYH2UOIlLnMkB8d0FuvMWpmgMfumX
iqK8Ijl5m7BNBVzcP8AWM7nW5sm46uzYlw32Cp5qaDtk+VTrlBwk3h02r9MroYJAQeKaKnnr7quC
SW+WImqUK696+mFiSajIoDIo1BpmOaR3Ag87dvInrmYVEqelW9RAMDC6wcXWD2JiJ25wcBDGueMD
OHDB8tdRFS9yJrOXCpC6ZphPtKesNMPzbf5W95s2lUh8N9GwMxqNyzQ2xJiedsqA5xnop+Vx4JW2
ymZMpUL6iR4po5GNenV+u2eS0aAt6qB5GZdyej884p24vgJHrMBe31hLGTGfgybQRPqX9hgZXFVp
eODUOizjNpkyhQ+TW1iKV0Kf/hYuyaifOS915jthrCXf7XSQaCOgP4+S1xremIO3PUyy37yYupOp
OqHIbNKEGJ8j6i4jsdMvxalUM14/7soQN2vh5Pyiq5Q18JxZDwOkbQi9m/PHKbF28Vd9jSVrwrdv
NoF+ope0iwUJ8ppiT5dnkCGDOFFs0wRwlfcj9oDsh7qq5cCWPxFeHaUYZdr+f6AdvowgkCnKxccs
L5puCk/aifakLhw/G9q/FW28aL2rujcEwn+Kvrgy0disGvaJ+Xl87IPobXvnZkPakWT8xS7SCluw
OAe/Jxhiwt9NRtrJBbdblSSJPiyuLc3w+0Wqt74LayQRKTZ67VU5dEn2q8rK67rTfP8h6uDLRhrg
dcoCRc+yES8bE44Abo83Psp2t+67g8TJ3ruJKq2JoveFFyEors4ma2bPZBkvuwF1NOVmD1OxrjWE
coVR8TmujvZ3jgLdR8Dc+YwEK/FEhLGp4CtjQX1a43a23QghpIYvjoC5K3cfZyPePYnQfHYMlXsB
yLfX1qjJuatd+255dL76y21cVoqTOQcufnaE0AexDVaqlYVbrCPtyHeN9C+JKAmBVkj3etH7yw6e
ghKwa8Hv2XgC/jxCWyCaKROidSy5hJZ8uyEMK7I8fNm/hUXs4w8Vuxz86X/Cisu1shuQDUwz2bJa
aUxU7dv9GulGmfjlQMvTpL0SCiUyA6wYe9akta4UAsU+jSJ+Eu8/mV2dvUonjwvPXPe2jyuAwX2/
8Eg+J3qawqZphicyKWc17hM67BZ0smhzvgXG7wQIphS/dhky8UtEUhm3hT43lCyc5oVhy2LhJi1j
LjgUeR3SSgBqaQctiIKJEOb+xWrMCB0iWa+ovDiAu1pRPJwmkhkPe5g0XwngGysSzxo5JbLR4ZCI
seH6+MKNm2xQlWs78+wpf1BkjtkBz9itZtZg9tZd0uwKlyEV1UOBnZ9St5aDzrJ7zPmPSfgdqlMu
QE1bWJbeFzXqblQsX5vSaCW2khWJX2unjXoqEURGv0WHSFZK8O5MWxcMYqsKn4Fn4KxA9m5495cm
GOrwd4W5DrVSsWw5F7j8Qh5+wkQRT1BC7sak8hIL9v/+g8uPMuYPmrL0/TO0IXEIbxTSR7OmYu7T
CpyvOLDzF/2AwrSkapc5B7AdRXLR0jTXE2wwIJJnQPS9lWkjYUhDaY64Dr3dO/XeSrked2Cq5CET
YegECRBWPCb7Hx+4+f/l/dS697PYM1A3g0VPDf0TjZuXq+HLxHcHJs8IfqATMryTxSkzpxTIOYgN
PspLXkrOWJ7uJcIqSIhGPNVlR/PQphW60t0JdPVa+TJuZARs6aaQeRbC19SAYD3DyLX09vfTyDUx
sUIC+NCwE4fjPYEeb0enR4XGRbn7kQ0ldmzTyH/5e9+cfu0QBMcUTn3ndDMvn4AeXRkPmSZGBoor
JRB1vOZWyqnozlhuzDFqZzW0v1kZa+nBYbwlaO2y72mLF5DZGtjm4aLgWcOtBOOtGE5fMhrPQoEm
tPiKCUGJnKzPzJvHu7AVvBt4l0IooLF++F8veR/qB7xjlJUpThRH3z6gIjybTnBEZ664Dh96TxRq
5UA8Ur9oafhcC+tB6wOrc0FHl6K5IUbRtcJfmDeFbBRxc0DcVqstHfEKEXRgaoOse2uG4RQdgdvN
QuU0q7K8hlBU2dWBYb6h/jEpQUHPy5J4Wwun8C8U4/hMgyuMFf6jJa3TCfr8LGyON8prIahKEQuj
7z3zo7zhkaapFz7nKE1Dc3cH9WnsfXHdw9Lggt5MvVeuECmVrRVer/8rL/OjC2NTXUYROp7/u5+d
WuNE4JnAahh33FwlNo3so/MZREXnmFrScQBAyTmBtrF2/BdZoANXVsohKLSY1Ltkhl1p17hykT/I
HIIKnBo603m+qTJ70yvk7WV1RYkb4tnHDLlOoyzQwGg4AiB8XvFUJUDhW50HeOIC2jHhWYcXcb4Q
oAMjn3MsJ2XI1hQ7byv4ijveurUw1sQraQJF7aZqs36ZYLWM/rGC2a4tLMTIYL/AaakVgQkKl/1G
Yk866ktZDO99n6eRF7q3C+30npgxdGUv6rahJSMOxVRR71ll5KqHpvsGDm6CNqpJhf6fvkYY0KAP
zlodW0G152p8sBawPRcPQ9dFbP9nKHUl7f9eUc33Z1zdL5/6uzJUW+9gioWtfMqpI5KU9I7l75v+
UOrLiEOksFUQSb3kZl1Ir+OopGf41ptmPZ0nvN+OF/yotgXiJV/ql1Pbpk6fVIixZOisL9bR1s03
9Fk8nU9pEXq6esMoW2g6RmTM2XthytvliztkVb5Xwu+TEmkGzzqoA6ZZcKSEKZswtMmwH0ljL8I8
JDPHTdNSulbX+cGaECMfZ2SztFcHfEWHFGSRe/YjUYJQ7SereFxZMfdpUCvit1XmylhMl1/QbNSW
yjKqW13/t8BvyIM6GoJDAMJ5NmsVxmiTg+Q0wfP2KflKTOli2hYt4D2phWrObpiQqMrsXA21R10Y
N8+9N4ck3LRC9XcaVRGWKNpF8nO3VFc/OpVJSOEyWf6DwEow9yfmOm/WcU/LOSJSEtVznaSgfIqf
umIzmpaC4BGM+bWxLGu+4x3fsKi0J5Mehhu1fQG1mqKwPM2I0HmglCikCFh9DM6rDimrmMUoEh/L
lbfZDm3SmkFU1xoJ/hLeyQtmtTNn0BSu7gNmaZwnLMtBO95o7f2FofFZecGSsMtQeQDnX3GURL0i
j8yXXVmTZneHMMsSCHKzIzVxx00zNlgXN0GxUIZRYcapfRgTWOBcl9ZTittOwcaexlNgLJ+mIpOm
4w9ZCY2+bVZlenWPspRSWcfgQZfWJyrjozZjRJZaswE6ea8BZhWBquBf8N+UVZQILEx+MyH/SpdI
yH/hSExdkDHvE6GXXm0SjG0DK6XoAkz7+y+xGMz5QAMespF22oGWELZavFuHqcjunQ0OnIk+Is89
xU432qKdaHTnhmagFJuou7nvW7X/Y9xkLkfLbs2i9csNuLDhPEw9O5LomODOYQTmV1odGRQ6wa+0
3W5qnZsEV+QE0iGsMuhuTKD8+bTLii4FTiglnM83s7hnvKG9VU76qB6gSMAIYMV4VKhhnUiaaUM+
3JBd2smZVu4wWflcGUQj5focZx1AcXjNK+mj1f6RKRXJHtw84jBDhIf25Pt/wpnWQgRVzEX+2v3i
RFyXTmMpraf708Bwhm5o+Dj0y0FWeK3zpbl7Rp+MBQh8GgRlUQt3wU7bevTJPjmsloZQsu7I2ASd
ZuJV2umLi7PdnW1LrdT4e5UfBY0anbjFXqOSTR1l1MB1ZW8fyMz99pyl6hUuh+oh9TDhUMQXtxCh
F3ZgMP/zWuyLZyxs7dmikZNhNoPIkJWHqNL2uMOLaag/0/otKMq7z7/mCwPMN8DhXtVeNK+Depxo
RnZVVkJ80pgJwB9AJAvUEziF7OJGx95N9fS8g2NJ7qJzkEzM3ucwJDUL0P4lbtwljbm8fibPHQNI
isYiyLClPuuOhrEFbyDdGzAvWt+yemRpXk5Lt+yVHbus53m51Hdjy6xCyZemOJvY1SY2ST869rBr
pKHgjt5VDwPvhm2VFjAnVzW4o6vIIZscBsgBazkdx27l+Pu19l2e987Zr5okQ8hR+l4lfqyQtFpb
a6ietlva4KvsVF3fKjOKD+11VBL92uahgwIQB9nTk56ozEoD7ljj7hfA/AOqkYzn11dlRrVeEqPR
PD2oUIEqA6iJXNczD0lhGT+1/rkw9EdURenoqeVkrcNcA+Yr9SfHzXXGgpztb8KRQJ050levoo8I
fK9c6kI3C8kU+9ymFsTtpF9pIC6hxiXLO/VgSMr6IryqKqCUsU2pdQ1phsi7SqaKKDteNdd3cT7V
HX/EsyGbcZULkhPdGizZiIcjLZa/R7cRA1+/mVzY0qWTdY2p4q6wryTNdkE5v88KR+HzpEnednpw
NY/C+i5/OcOJcf1o9qNa1cEow47K6vfyx7kKnaY+mxDP9HkAaRK9KE0fWBAimaK5LE7gQFIsiCPO
L+b6Lw0P1hQudLBmQSzk1BmoSjKvZT4zB8RacyRfePhbOrXQ9e489/JnosLkgOkjapuDSmXtMJYi
SDu/jGWtuwUzQ/cGDj+CqozCFRXZUmPcYnAdghZ6nAqFFQ95tviwnkRAFpkJjKqqkikKKaZClNfg
QHKbe54SA3yHU+ZseuQ+j4l5eWxnVBSYejQg98J0M+CoBMGxCZlJjt3fdJg3F3epvpPivXJ391ns
QzOyigunCw+ijgBfgBOTzvKxR7NRB9B/XTo+eANlqwU9ElOq1VUXRcd7RjnZ6siI/4/ButlXQncu
jrimrl0V3fR+IutZCJWqxzpXFiNd5AzzVhGpaTM9jXX0Dg1/E5DyxrZDOZ+eBDgYrGpzgJc4PgRU
X6Ac71wqdrjTabnZzZRecpU9WMz/OU5s22wHxUtHHjaUJq/iwQ8+QYNwVb5etiSB9bQA8SRcr3fk
3LFbjdjQVcNc1SmGAhHYFioAI5TmRN+4ljZWvxwqeWW1yqzWPK7VCZHKEuNSKbr33bAdZE9WcXkU
G6qyfs7HYNYG9zGLrRdHuu7iSI+c4wYXnnR1bDCWFabkd/EBketeJJTs4EAXu6FMSFjNNqTz0P6S
1hqIdUnqJSMiXXYVekPhiNWJp+oPWLLijIVLlAMC17BMboAnCGIZSonptVNT8Xq+WwbjZWC/JT9U
mx7/eZUlFybwDm8QVB6Hk2i4CsDfEqxxgD3P3smVLrx8V/w52PV5xOpDTYhUrRgi8MSPitJ9f9vg
CFsYL+7ZL9Ngsj7ubdfn+kzj332+7Qsje3wkouKA2yw6NTYPjlOK0Gm4QSYEGGN1xWRQy4eSrRRu
6zaGHQVEhn+kVWnap22l7zSj6XxOGU47/SyUlWFtmJ7E/39F3bmDKMsbBsf37CDUHFZgdnsxLdVx
NhOcaBZgTuX6dB7U0RurCMb4D1WIMYqYoh8/1nEh6rjO6lJkOlAT4G8ru7PkYFSvE9Itqhgm+l7a
Mq+xsXrGk/YMfyaKHVMC/cTFtvbMtlCGNN0eZ9cP5umwgp9b6LsQ46epk7eMKYjxrrZVeRPgzDvG
7vYU9mVaSswQ0KV+1fGOCfK4umk/AujUlChapd5e75ZCgTUeTBHidibFDMmDHuba2mEL+SX+a01X
uCRrMo714tyj4xygQmUJVGGvMxBVDYiKTOSmuCelmEhYfNHvCG0NYnjBWszgr0OpvNR6WE4EUjVO
6t1y7mrCgU0G4QeRx8+JaxmQIV+QWh/dHr51gRjF90opX6W5VyBp4bODM+SG1kbwKFi1q2zhLWsS
eoSGt+lCHaLv9NWfYsFwKvwcwN8a43QcKDEyQuzKQj89ovkNy5yCpFZPUFgrznL7fcxdK8HgOlBf
xJIrwqoVVoTg0zrIn95lUCqFY2ey1TNHQ1vTYu7vSDNhZGzXOiI3a89K6kfC9SRRTqkhYnoHcidi
ysD40tFiJhKO8y4+rf3pdQVTDVwCGABK58naeH9urKnXdV61ouXl1OXDNJjYTCkbfo3DFr3/JgbZ
W/7QehCd/6gZlVe32amATV0deUfWBNGVKvV5Izg/jBiFAHLloxy58LOeZH+czeZET4iAgIN1UDKG
mizvJf+ihqapp5sZPuv/fiOCBkNX9/iFJnxMYKwegnzN6IJ04CPliV1gm4QCWffFO0YCPjSJH9cL
y9pmYIw+d8Z8UaQRmwgQ7iSNTFfGlbPTxFHlfG+wU2G8Jt+s0ypY2nS5TlH/XwQG3Ce7LiN+QE2Z
UsQlM2t4jEDUEO4326/5uxSbBQ1bmPUsym+2lFvMmNn9TvAobPRd0QnzrOAtz/xKLkHc5DMKtXgs
0ieg3FvyNwLbJNriQFUwq0pQAMagUtn5CzeLzf4QX4KZ6QvoT40vXZ8QEh1RhA78XPkKP3yetZSe
N5WrgATKX327qPl7JD6Wp1Guk0Vj4eURptSBqOHsJiWMW0gzEkwH5t++ZIQdM1KULpHGnfG2vt1c
MeTI48Ivz9xEQRa+byV6nkcsXKVI0+uzmBdOwhvThu2Qp59YykCzfqrhdbcLwqFCnW+Jh0rGqj+D
bZOOhiwWJfeE08HE+rvI6LAiFX+Md8Tmq8n9WaeNrVEdDQl+gGCxiiu/cX8sUEaq9knRRrXP/dwR
Dx7dGfmjujJ7vgP6gDk49FTuf3lkiAC21UXQcW+gyfFQXio1wYSMQ8eTqygYbkR0nbuIitRpgeqF
DLiiBa0Oe9s4NkA1WYk2RkedgYRcs7bRhv0DNMhlUph+VtXGWPqtt5Sl0iVB4pzYTwxwW1Gdlhfk
61f5w4g3YpvW+geBpS5XmgfzUNhz2uxuWtAA4YQZXLGXalC9gGFcXclxmloN3g6qLQavo1jhh1s8
x6TYuH24hCUpVAOCIpnK8j5Wfum5VglnJ7Tq25iN7jvd45SupXxOojqeIVIqRzepCjP9bO+EQ4jZ
3sh2bPlLYi0NG5gQtI0Vzvhx/i47tPisWY6JYYlBnCWeaY3WfVjPtcwyCUYI9/VYs0/rFk/nV3sk
qxhpFKQSAtZP7+p7Rgg5e9V/MP7YhrcQWhQJ383r5JwE1aNs19aKJnv7GwbqLu7CZnWrCO1BoMO8
7ffdxKI7NvS02SXPgWrBX0+rzUC99HBpVn9n9xTvlxAfE8GndlBIIDmFtaqRTBdYFvw01Xri13kT
FRJ2g5j1a2CHtxsO6cJm/R2I9cW1S6WWgjxkFJe8ab2dntg2RJ4FOE03FgMJl6lj3ZkYns+hUtV9
jd6iQ+1V21fUAVDXtn0/pYOfWI/FRCNVMMhJFn/FRsmGByfejcmUfKZm7lssaRWk5lsEwqFuHf4D
7oEDZilvY/1/5E+Xx6uEai80tiUvmnTWzZzf1LMSk9XmipezSxRCgcHDjGHB3PzBcIFeQ7wtQZQ/
X+LV5Cmjnx6wCGAbh5cihAKHLkneI3CrdWGB8zcXPunrHUSBl++DPLDfg9WKLUkyOqRqITrvMNh+
SSQ4qorzzEad96WbuRpXcRRchwdZ/kZyqSLKxxNr0YzTjZRsjTH4ictJwmCvwuwv78o95trSM0/W
Wyfreaz+Oim6oju0TJUaDrRPRUZelHlCPJECTM6lhQWry1NVGJbAe4m2BkpCXvz2WD9HMVowJo5x
Rca8t9Tre0Bvru6PDuhng8bwbtdhzXtfo/zxJFMYK+HNbrZN/jSHw3hNFds5CnQ2E3Pchj3m6bxG
26gh+Wsl6ElCQR3ZLdZ5wMstaeSqljPFuFB0L6PyULDhswsRNXstipnGP0ADkQ1D++cVzLdi9Af0
fuP4NAhJXR+VkAgYAErXSVmLdID8RmftydXYoSYTQ1ArXsZzwM/e0jzyehQ4hjRResplcqmkvKjf
E5qYUryINHFCJbp9yfa8YIXLhyVpqGi2kYTYHeZ81w+sZdKK9lRJAdump+G1p2Knyu2m1i0bDuEN
afBlDb140peQ4sJozbJw5I+ZtTD5mKEdYJwHENQNsZf3nppihmzubRbqsuARFcqu91G2V0Ak83Hl
A+hpXUJztoK4ProlJARRMsuldvbqvfvmgjAGFfsd16J7gLX6ckAT1+VA7zZxjxlnyS0r2j+McSEr
7qauV5qdsdamf5Twx67zwo9dJ0g1fV792Vl20B9AyVR62pkLOcDBlLb8921qXKocTvmpp1wmCT2g
u5xiufSDOjhEtqD3dCcGkGzGcgayqEQAB/esrbtkiZuS7OH76OaqKekfNMVKALy2R/KKCaTiRB6G
HrmlarGAUyhrxttAZ2l9L1WExW1wf5/Q3VJPXr3qz/by1iSwpaZC9c4YD5laukgrSHzd5CLpT0bA
w9A6oBNI/vxBdQoLPhJE3GwHyjNTnRA9V5MzTg+2wemMECsQ04h99tuZZYa6qo5JZoWRL7mKNizA
/uertTM+FLGi4f9vijIZyiotw1ObipMu3OcTfuRoJDjZi2F+c2hNHs5wyLRCz3PtxB8Hgit/W2Nc
yh3Z8ojbgQdjJpBNZhXz+OR9Rx1EzM4EvQZ0vGczPorG2xKcB0s+tKq2uGlevShr6mfdDkk9oj76
Ri/XRqmkh9I0AlxhpTXMxvsy1+0kmGdVb3ZFa591F9Nm+FqSq5rpmd4puDg0WwOSQOQiCXS/3iOf
fJ63SphtsJw9z4CHVH6c8JFwjdVgiV/uEm0zPYhXHLsY9/IXqwLsZrq6Y8HUr7m+F5prl812j9Ag
gSNridNnoeo+KYYFh25aiNSs+Wjz/5W0q9TTdYbAHVja7G2yV2Hsl769rBrcdbAgvOTKpLKIOz5J
i1+z33A8+8byNnU0aeG8YS9H17CLd1/Gyy8Fvcz3zz/B6ioWAnwYrInfIYIXzKU7ezNfIIquJLDK
vZ5PLndssrQPiYiqKus/bsuYnNld+u9mAmgFMXq7l159HJ8/yeyunA4Zu8YUvV7usJfueWf19H9W
aVpSiQ1GYcMrwSIuoZZaTNHQNFj7WopK6JroMN0AgxqGf0l868cRD/ww9MjRrc+SFheJuc6H2wpB
HR84WqzDQFA3w88FL3xFe6VjJ9Q3zwqtH7azzrf4l1ql4xcDJj9e6MLVO+Kbj60I9HXYUTRf56CB
WhBmcjfa+Gy1sXqAVv2+3ruwx41LLJiKgUk6DCkiZ6ZSvDgn0kY5btzwaR8YsY2twFRtjvhAGW+i
3VQTcDqd4EUuH4+vz8wmkHABCoXChkGbMYtmkENvJs+sS3nI1sSVyi33duqaHpwOmzHloYVq1UAy
osdbxm3GrwC7hvmlqS0MdRQ/JWnx9Wvs2JA6jDDbyrLXSUhe4gHxnsZhcX6hl+zGzUKBuiErkmMg
BTItXYpt589RJWcERJ6P4r8HnAMlY+fFqdTpcxSnqUzCHdJdQU6lA2vqOVd7GcRarnA7iQsxr1LX
W2l+GEU10LqfCD5lSgStpRxLUbmAYER3U7kC3iflXwPuyeptGUPe0/Bax2bkESNwQEnbXcWPvU4g
oC3Xdci1Fs1mQFPtRh7wmk9eKhrFL9AjW3keedSyvrYgmZeqDZtmKjT++SrUsl7EMqTkVPmRz7lA
H31vyvELsl3BUqxDzYau5K4EbNmq6XNj60wT+WqdDlBuDRU+pDf5OuFjwaW2WloXrhk7Fz4kP9ct
GmrmybVNyPoyGFBCfXySe6OMcNTIzEFjdaxGZAZL+eWKE3zS5IamEsTjL6lQDvMsVOP46D8eIPc+
SssFJjG7JP6UaIyXb66+grE5Wb6VehXUYTycsf0hYqTzAeUIWqHoTm1uc1XR4+3raJ/e/obwQDaM
TMvwyG0jP9j4iFCdrqWKKxnFQ0CoLeNiXdKxvF7GQQ3LiVePpdfShZL0lcaLyYKKpqFd2BfH1CVS
hA8cJrW9sdo3U7qOY+mTBNC/K4TFEkOKVY6otz7uhU3c2Madau6A3+O3JkxCQT40irGOLMXwJUq3
wnFfsshZ1JyTUNGkLYndVq7m8HbMRfbv1+hQ7s23dbM1FOH8Jp92wKK6hEyjqguMyn7XogS6mHgr
7PxfC36Yrz2utiBq2QiHuoLflj4get5WeMKaO4dELhorsrNIoA4NDzF0Jp0iG0iaTShfRhig0fp5
c42dXbgf/faOX/gICozOgmhD1US4j2N9MP/0XBMWAP7YuCQVb1S0KhEQzvprY4nyKPaKsvtSJ7aO
8vD8Qy64GNaRhBAPWnuV8LQkTe0QY5aLCnGFFvTcI8YAuBQeTsLdDVbVnIGD9mR8RwdQmcIIQxVf
JVse6+LExgYdcnaSKYcCzXKM9ZZxzW+NoUwAFfn1/puBZQe3i1j8VZeXLXkerpGa1V2YNLPxC71r
7txuNPS5EwaExC6oQHNsdgTpuP3uddkcfeFlAdLlGsmZ1J9N1+vZlET0T9dg0TdI+mFRsNcZwhan
YblxE/WdMniHhj5zxbBifqxoREv20TJDB+B/xHUWCZqZ5ogPzjAASAq4cpMQpk2aFV8xf9C1Ps8q
IMpABFsxWvpggt3bGIISc023XDaAXB91EFFOSGHS3Z1xkHpw4LLRpXPIRm6VJ4iUzidt/zskahQt
/ORSKSgDBCO3Y0m0Nhlj/XvE4qYR+I69AYc0v97vRPQNQnxfyiTq5e6pPUwsl9p151pugxrzTBcs
bEHM+GAlqPP2ecGUJR0F8bnzKC9NGWwU+Th2cN0GU1z2M7EqTah0c2WJ4QiPP0zMZoNNioFx39iC
XndZOB5PeqoA887L2CjfTD7rVFxC1VFkw+JzDFFzo7f10mAy5+inMdIAhweHxxkeupThqlPn8OLr
ym/CLfj8tx2D2XM4AtddJaTrp8AzFiSZ/lMYtHsG0GiF3f9btaw5Xme4VVgDKtQUZLcmkXDV9p32
jzup1iP2Z/hIKzvrvJ4Qk7DniEKEiI6hoqSrZcx11Wnv323ZbTyx/cI5RfNyVGSEyxcJ/X4e7aGD
FPGHkEx4ahvj8egpeJbvnsn9Kex9JkPCVw8BjUta0YwzPG9AxaPDDCRAKpdSH1P1xEcdKLJZcj5B
RfT6ZA1FbGGNI62ODhdAwW84FAwuLrLuMlg2tc4UWOvCdkI8baMvm3NQAODv1ziL8UFkFInfUHef
hfo8bRhh0B+TkvR4ea7UoHbEwkfbGhf0GIwSdnWNiiWaU1V3cKaCUzSbO08GOxAr20lL7r1NsjHH
Pm9yk+hsmb335RHX+cCoXomAMHTPVd/3znRsPQXBdLUDUlP6QEeGCRnUHvdySh4hDJ8XKICag2Kv
nnxGCSeiSj/Rc3vxDcyDnaAniPduxxZHX9Ig0nGERVph7ttReRUpZ3oYb83A4x42Fb1sc2LiYqDz
edv1cZ/v2kW8NonD5zqiQuxkCTsMxdasmF/DnySNJx7NtL7K6OYbPsMz+uiYWesXSgLaiSns2Dnl
vlzaIOdMZydCUpnaaJEuTzGdnQxRLC1GbK0FYl7Wpaym8xU5qkSpriUGyXSQHfY7I+Zc62nnTcT7
7DcqxdYKFyMTQ56/q/SAiPeA/Wv3pKXmgtWeYpwuAPyiwaqWSJv5oAWTKrp4UeKFXgJU1SvnVMMj
RL+YcMO5VtMtI4OlrRcBKwwUG3ZjREbyKmk54Puf8Cnw2/leCN7Y8+WgofIbptVQdlMqGwBY2rdx
YxLJOYEcisjjyr2EVXBFSX8zwkxqCN87z4LgcjaT4BsEdHLtQdf1lhzgYswrnlQvXZfQPoV3aJjh
f0o0ZxAkwqaoQbYXH7jL6g1fYxmKkx8Z4DtlFGUGY/yI/rpjlglrgy056NMQHww0tvZRHhxfY1sF
aw6QeMFefh+6O+g76xzBah8ryQWu84Ul0nuaDnzjEdKQ855UdDdRiw24+WETwGRNoIA4V8qw1mqz
/rKj/TaxFodRI3deFZlfA5pJdWaLh4cQQj/d8xlIvWnKU7trrsaqrLS40t7WeLQTHdBGOGhBoPzP
WWoD7WPBN4H5CBXq5AhBZRg7/1wqRyGReVQiN3g6MUOXc9qkDlkyFGc8Iv6AnsUvFF+n7lqArfRc
fTMVXzPyNH/TPDie1E5FjzXk129KY7rrl0ThGH0GPpTg2jn5Vx30dPhcc4NNfifMIALnO+xyQOdb
9bMbIDAbVGqxs4aVESZdJCMSK34taujRcj/mrpr+jsSzy24CY9Xi7eK4LZtwE5sVLGPUeWKY73rd
ZQ/jNLB+Mo2fHxBIKi/K1RLdJHdYm1BO1cH4hjsnHUkwv/sMtv6NlcTS1UWj+O8l7b5MkAUle8bU
OYJJTRdWYUr24teGmYcS1Cv56lJ5qvZffn4tleUVKXCczy4id8rVnzo/SL/qkbTZ4OaLySQjj8Mv
5Q/5/vGbpWFBHyIqJYfx2HHEB9Y0GjyONGTIDmrQf1jaYucHS5/n4WLXkJu0rXd4xCB/81oMriqn
0MhdXksZghkzbRsLo+tD94O+pGxrrqyoQvEiPmdfl6AJMrnXNCiXCd35/+KElyF2isWjKc/fR2xb
B6hUi2XiH/lWyg0Ff+zAP+iqnJwYiWHunOcHvS7KMlbxLwWCAbFOKlAR9XYEMtXoge5pkceFJL9S
+3cFbMFHUDZIpFTJVB9PuRX9BU7e4NE0KZmMHEYEUtZKzOHMyTQ4xum3IDzNlw2iJqHv6dt/Xs6F
tQh/2ZZYpDWyPj6p2/jCxZ9bmhK7kqRB8J/G9HacoXpFgXKL8T4h2KIwo9YIamL4n1aHrTtZGGf+
jV17IJ8tGjYovQNPfaCXAWodjbvwuPYH2X/jKGbGyPM/JRZUD/u+DQXdP3PCYOG+sSq593Vn4Aww
6aTNuG2W9G04uytIxWW/dH2tuMMtX5N5Bf/ynhXHgOHQFjjPVqxr78TzTZLuDjIWC9xSY7MOsrRg
wMgX7BzzjTykMp/+ptLF8W771nQHN77cAIUfQmI+qMvn91Yk0xcnt1Fsme8E/M8t46E7TGqXTWEF
mI4emLkiJaX6tTvs2QstcHZSGqx76DbYoGvXcUG1+pdZBzdi6xJnj1Dj5rJrH23/yrXOOz3JpTml
u7zAUTjOsuIy25JYDE1KfBqVG33Oxk2bcbZbf8LvDIkXDyQU/e0aObVxWhfLfDiiiL8uGyC3FLBT
cpCcIJ60/5ROGHOawCTbNqFqw+P6PfLaLSZL9ro/hjXTfdMY4/JrhiDLRgiMfIe05daD6RToOGc0
+wCtQ/F4kcjxUaf0smuyU3P2QaPQmo8mUS/bIkVUDBwcGsmKM46hLRbF/zeywH8R+NgvPWz5BkrJ
9UrFv59TME/kmjG9sNJCVwkYsM6doxlTLgx2J2FIP4EW1lFulaDroxGApKfALxkoDKk9rXW7r2ae
Z/jWOhjhPuUf75Wi17eAFMsZs+8XGEWnrSvXqCo3GZyiUr5b7V0d9o9RMJHPHDPc74Ex22JzNj1g
3Gf7IpiBfzfcQODhUThLiGoCoRWIchfdrbE9O5PkOngvpqqmV5tQo2POl7sZVA89m6bVRNaS5DqT
miO5sphoRjhWc0MiyuUcuTILfXc5prWX1s+2y3duZS8btBbHRPs6hopgRZIX9fLH6VPWKDYf2Yws
lJR3dXweKYVhCXd69SALvnSdsUpvY/h4YkWJy/Z40xYbd1sP0UfgBslA2ex1dcIICNpCnRZq+N4V
/4cDnbzAnCe3TnpgFUoOyqyBkANIfieHBr0Dp2FbxA698XA5dPc8LzfSm4nQDH2smQQ8L08pmxAE
S1j6znpuiYlxFiE5/gTeqCr2H1IG/xZkDaX6Pqnbe2FXFu0CyA8D6v0GIcbrn3KfSWdv8b/8qbTQ
9DBPxZ06RUeKXF1heeRPxF8z+/la3sy/HF7+dpvneio1XOi51gagci0jc4LaSoRPXqxnStaRoAV0
0Be/Y5/ruBUAH29qr/6aXJZGjlYmdh4crQtMvkNbrNNIQMyIvDQqrxhZl9TPY5wp/jmGVRKQW3pB
nfzgLXu57YOoKc0OONKXz9BBJ9Gv+mLzAyhAfbvojypsiPTg5j6TpvCLmPw592QVOADDRHHGbJHI
YpPbaoV06S2o3L/6pl+neO3N+lGIZ/axxZ1sn3L/IYLhKGhgAGpuF5DLQ333zqXfPiUfXP46JyGd
VLV9G5T4S7aMSSptGjgEkt2KvU/azwBYiLw+IOv9T0sLKrWzyL1tcxoFr2P+NM95jvyElqM3x93t
GXpfKyBKQU2K3jSpEQ9zeKCMxg01CYX/NMYRrrvMO81WzeTh+8xxO0tcYy13vjLqt+WjQb/b9Nvh
t4Py82wrR0rBQbw5+nwsbJMJsOHv/8KZ6onoL5hku1skq0fhxQ3Fsv7/kf7P+FvqLcqcsvybEgli
e7KKv+YXlmg1g97197HTzV9M+9xyC6LNWh88XPRUMH83swoQ4i2fepCSVTpeTiaHSB2hn3ZazBZU
tHfvwjCGaSDStHVMx2tXxZW2s+Fu633iLtLeRCgKd+mAdC0jE48TRPP75HkH1NXxsoa6Hu7j7nRP
GFdcJy9sBlYtZOd0HnP56NxVpSDRmg6G3rMWrDBhb+hGSzDRokG48NTwLmWRuJ9eh3NlsL0DA416
LVRNCVRzKqO7iCr1AbrfNimds+jHU89VouZDPTqa+BQUmKVM0w6+B3Vl2DzXpwrjxNs/oVvgVom9
DTTwWCAo25x6L7jZrP8Lxu8i6jzm+wYykbZMTESwFi8PErRbkx0yRg/bOLAP+2auvX37Vl8Uz+Xt
NfhuZWT25sE5V4vlWccF5Q9FQCCCEXqGmxvMDuhEDsXfzIcRMuWqYUNF0JleG2J5FbbnH+UbCapA
Noyv2I0Q8jesTSwIhTC1+P1Dc6mvwZgS813psgiMbaChq8XcapHbUGfJ3rYDcWVrY+R2GuOIth3r
ja0WT9ScPo8y1SyHP7/cuIKqZ/WaafXDPa4ML7LHbPE4phdS41/ySO9P49VWJZ5tjvLZ0p0xnjJi
IETJjW/G1DXzww0O8QQF6qomDL6d+gwWT7VGhlcF7DgiYIWRAEx2bp0FitataJmDGBEwUyB90gNX
e736yJ3QSka2WeEL/lPpCwdUHv9GMUcgH4O01QTyfZscUfX45lKwiZzCmL9dHUHjWBMJOC5RIjTj
ay8Ir7aoCCjMfxEibHthk0wol0AYtEBkj+L7uppGuTJzd5ULUCzYWJIMkAYHLSBsp+7uTbXBY8h2
AFEJPedkXwYsse/vCW/q7oh/bUKnRrGfP6WQtI7LSug3S1p/++R4jibxT2azR9KKicoqnetaT+Tj
EFfDo4OqPb0Nzevm85UnTUngLXwCaLbT3hCKHpUSqpDeSk5j/kQZYpNNi30UMw00iIGUNFg1cB6G
45g45LqXnUBsk0/AvlX10pXJYB8LWUOc0TzZaaMrb9jzzFvd6kSnr7Ew1bwWPEVRB1SwhR+F/Hq6
dC0kKxO26AI8Zrzailowx0nW+8+rZcRtvc1RtkbxobGeov/RldzJ3T/FRp8rXrj5KTicD37pB/iw
gVsHwmEjBObU4GVFoaP2NSPynkM4aOTPEUWCSjZHKasUEXQXS6vDu+3drMzwqGZF5hX6QcrbKInF
7kWipEETBTJj476qJTI5yKUwlR4ZFffzZutSfhen5yLxMVRTs5znC2IjHKjw59ahYuLLvGTovf6N
ri3TnmUuLfx01ZCfABu/Th+/Ri32tQTy4KMURVIToraTtexsw+7KlOdExuX4AGO3yh1BVerAciI+
+o3agHe/fR0vbIggxiqlP+KfgJ0QbcsjrpP2gzMnnkDckANsi7FioWcxPcdWYf/IMvcnFlfrv3il
SK68KvfeTnUCWBVuuI0LSQxl/UJgieconZsE8YhI9BsAbIpjtm7dtwxg1rJiB6sCRFrLJwVKL+//
lhAq+Vn48P3UYgzo3Sw0NirrnazIq7DnsWBD78NJZwkkoVfeS+8ihv9iYliocVff8sQb8gEBIULh
Mr3e4w3iqssTsfNeuseIHZODquP8dGTzO1wzLVhN5aPI2ToJcfaJPxKyFis5pxSstBfCfmxQD57X
xWOogt8p4ndUmeQ/FQ0fJyE4xle4ynZ1ZsClmJUfm9nC5B5QtLcMDiivzeknNV12frRkE0VpiSVY
w3yF2pOTg4fi87L35+vg4DNNx+7ExVOKB22Ywj8jK+/vXKr1n8EUaOaB+9i6WYNf3YZG76HnBP3v
DPAWmIFN5hst/nOb2/nPuI5vFKfc0TnjOSwz2NZJ0rfZewrCNju+uUCXln71r7X3bZJAFjmJmsy7
Talpd5Szkab1YkVjDUSlqM86i94RGprexxM9TnEi0R95yjP+LyeY92zKpdEXvUfhWNgdY8eIjJqB
G/ch3oup0/xC8jZx6Aee8AP3uxNtISTpRO8P06COfzskxtT3DgvyVOq0haLBnwHSG+kYYAJf2Wkp
CG5q6+lQ3UanSwK0JFYg30onhnrKTtK1Jg+IvsZEFPcSfIH7F2VIF8khx3eJ52fs4hNDUAOb8CoN
p+KyPTNI7ubSoyrLxCqs1NLcYujgRY3y9jO0W+6qpTpPUelSz6HgM7Iaqr+SuuEo6skP+21Fm9f8
ZadJxW0k3lTHII+23FTerMxJYCoe93M2m1UC+on2siWgK9gDNzwKfrEyD6CWwR57Mf0j2NfDgEjt
yG3jGKk51JzWMmGMwK+uvYbSnpuBIaTlwfJMXL0HtV88HjJogsOjHC+JiGBkpVpVHKzMDVqxSflM
eAEjvnLyYmUksu2Cm7KnmeWssMF1uslSR7orOAAaxPV8sj78kEShd8un2IDWDsMcYJsHgLI+7FC9
7L6nal8p58mqFYMZYTwB8jvASm3dQjLZKB2XJg2ZY5PkqHWiq8X1WM0tYTGpw+iNvSTMlBEXCk24
cRruozcNgufrxjjp5qnixwM/uTtdJshiangO86LlCkvuBe0hu+oXJoEdW5bBXWtEgQr3rFhUNNDx
UOtU5drbvDIicb0hfMtDvYVTnBigay4vzydZIq9bFAabm0Ppt+Ld8uk3o64LGVCqVvKKDIHBASgS
PdciDnpTkIJlqUjw63Fp6gkibIMhM4P+9lL4K2W4cXElPoSB4s0tA7rw/Hf0FxB/ZPDHL1+fwypY
s+ypHA/6iVuuYTqdH2d5+Zo277+X9o9xTub6sYaMaJ1rDrIDuHma5LDc96qyxbkJt6e1WdZP8bkn
B6HWiGSi4QMm3+uMtiYS4bcswlwWE9hXJmh4B06fsd9B2hRtw2qe/UWKQWednR/PekV1DQIeAo3N
19ONZgIMRvhpyZmT+FgnPzPRvuAZtvWsF4rwUnyub1616ywnP2FkElqc/ZIMn+jvYFDUjs4Cu3xn
esCdHgm8PztnpL07tArPOy/e8ig7RqoZZF2VlYWnIygl+RZ00biWxEL5UOVPRnLUgzZ0XoOLQOmn
UtihmcmK9vhVv0Rh9+8Iw32sXKtnBhQ+b12armacUqWjMeATe2vWNqqWj2nlW8Lg9YbYT/swZvPR
O4fJ+VEqbt9/XcB2oc6bZyeMkU8mlnjY7odM1KttMl655js2iL3VbK2sLb8TOUpVW+Wy1hc+aW+y
rWSlVk8FWWfcHycny30ndqrfybr2gmiPAuKG+oFphjEzFnMOGH5JUB++PLCGbksckpJ1nJ1MDEkU
OGIgTCsL9RI/nZosVKjMyYdAzxVDR0IDBg5zaVOF2DxWyu35WdvkOBGMmrr8DfompdGbbjKQ+iNX
Z6BXjOA8uxrh8MPdkGu3WugDKLyRilzIKdwh6rmD2kooo8DEcRY1H1sUOY5y2ufrWkTU8viReOYg
MBNz3mpqhY56WvbwG8zpXrfjjzASgH77FJRrr4I1ZNwUaOWZRPg/S6LgoekvLwaWkDbM7pKaeAlS
SbAi5ksq5mP6VcKbWfYwA8wAT8mXrwnzCeBxSpQMW66eeWwRuHEkSFGsZ/KcF3uu4sjBxybYcDIe
Ow853RAcq9qnvfTPxXkOPyblmi8F2r+QnpQ0pT5Jjr/w4TMK7AxgKO+H0Jj6mqVTMWxnjpuZQXde
EYqzzxeObO6iIWbs5MKcHi5rxJKj70FyEBuaJ3atdyIZHG8SHK/BdZ1uT9O+BH8A/DxvWvU516/x
XyuACHRZocvVyd49FxHTPgNe39Yb2wnQZkcE6ti4X36SY/FYC2bduo4isxZgBb2r59DPULSAwb3G
6VCOInG2lO04s0UyRVeBydRHe6aaOx+wuFi8vg5LuFtCvjSijN1S16fAKSwfA6plbq89J7qrOxWx
QgOwJlTj1/pO81IPJHebdCvpVNeKh1tMdM4xs7CNsGoXaZ0ib5HakSXNexq4a7HTeXqPas2XYlZF
w3L9Pb3epkBAZWzjs7WwlOYOZyUKlpvP8EwxDwBQFzHPDhUJLvqF/4W+nX0GaSF7GqHZGoTdSE3P
cDErN9tsZfxf7W5D9bR8I/G1PWkWA6Cgp6FHZUj7T9O1IsZHK8mPKDXRjFTPTgWOg1WgqWNkqeN4
UYPK8yqSo4DIUbaunzApyEbN427r1T/AsBrXtb0/ZIwjOrjoYvgf5OBi3XdveX/uR+vYKgJggRMX
9S5DYm9NIK5dY1IKjLZzhRbvmXRidyqbCJGZs+txx3L0m325F7es6P4tGjMnXTCPIyDwUZXUNnsV
LdvP4eGt63r8RTf41CbPpBwWbrZSw4a+6l8uRAnv9Zu9OPoQBRWHQ0I0htEF5Fyx52pHexCbRbS/
5G91Xnx/Lh8ZxMolz1dCZZUEOwJSfYMcb+iAtDMWNXDrz4cG89DCFSAGRxv/4we2GDjeCgZ4NhB+
uv7C5/ExYoHQDE3CBQeHmrEHuWB04HYnDTUsVgin4BLWERBit+96ZTEHMc/j6JQFq5ru0O8HUpf+
+f8cxNtMvxS5v+O2CxWUd5SKLTJrDhw6OfPIGqlwTFVoi7pL/ZKZiSMkt5ILRztuaym8tmiKQmSd
L5R0K4gwIUeiTn9oA+a/ew2mbSm07w68QayMqnGzvSH44+pmnOR5uovRgPG11BYTqd8lUupzcfgX
kN0mEqwPm+CrEdaJB7XT4V0tV3iC9RRjhiLLSwCBFCwoqseTk+LGPYGT2JKUM88T7yAoRNUh0F6z
E2Bz0JFfjYgrC/uUyzC/k7OMQzfziYyZWphsW1kpEZs7aGYKfWhK4xnjSgyTC4kvNZzjPpvJvTHe
cuFVLC1hlcZuccfmJuOl/Gpheoi15KD2vBi6O+1slQbnsxnKYE4Ppj1Jik/CJTywsZAlg5AWtjih
hW3eyQP0j32AT8ro3M0C9pOnfAmymgK/z9WAEKciUnhnfrH6q7CVzf+iVz3m0hhkIxUoMH7tMwfs
8H4N+yI/hZKVsdfzIOKp+3BYYGYee0zC/KYnpWqiRcVp1HzRFSLIz5yBC0MMtme3PZHHRV3J+CxZ
W+3RgN5aKapsFG+W3EaftxUAWUV0BrqZAoAryvX6+iKAFzyA/kOhthivrLrKSUyN5w9DQl9IG5UY
LC5anq2Utg7jMfojTRAam33hpBdiRB9sXyBqUISa6GA8TZZF1DabO8cRZCElTGod5TKzhxLtOFGK
RrNauCEgc74WJQyoLuw55MKdAMyn/PWViOtNEai0GCwqphL2Lb4ht0VVE7/YZpGzf4/HB2E3H1zE
Z973WD3ijiJPSA1Y3F1jA/rrPz00QgllZ8DHO0j2hpDfaKp24SeGUh+mPTHKSz4u7VKEKfxGtUsQ
MQSsJ6hYvDyQ4xvZ4YSmETX2mxtEcd5jkh3DQyhb6qvRYqPRtoVOZyxGyMsE3v/DytCiD+i4X62S
nS1/NPWEydPy3bdsmDjZh4Po57xJglsObQZ8JaR+MIrHm6BXSqiUQ/FJEaAx7uqRlxaQNKCa3EUA
hS3T7Qv7KwVSR/jjMPeXeh847QzAXkN91zpK2HBQz7DEbeulni5pPclkRhjl8VOHi0e3jjhEMd9V
pgaD+xRa31uu4teOxq6bUwjg0VLvyJPJbspKIJ6mNMmM5agNA2kRDmGMH1nYJyu7liV3m+lfEVpd
eUTV2OKNPnNvu0JXELzM0BRrA73oo7E6rIrXX4HqhfMbppPM6JYkaXMGT8wmvOsYhwYBAS1aXbHV
2oWMVyyaoZSP4HsbD8hF7P50ylMmByYRr5tf8Qhe+yaFB5lSB/fbbQrqTHbXHxZq3Zk9KY+pvImL
SyxevP4JrEsek7GPA5YTnsjj7xeGKPGq7ST9WNpAG3mCIbNqrP8jJPgfVouHGk9PGLnaDXmPHW+X
IpfM+eVmL5kYRIiVdfCIPHOsd49XirX2Pmz7VapFW1DF5B15Lkapf/nQibLteO1unMvm7LWxWtEH
4Z4T9KY0hytaSSzJKW3VqYt7NDNfPQ+elTncgkBBGIs522gxFubC2Z+XoJZ+/eZiFHF8WPNfR0gt
aHHMSnmFvnWGYlXKRWM2HJz4PMYRK//pPHgDPiK/qHyHMDhL3TGg2sJCof0kZ0qHR43Ir18a5a6q
gEUZ+K89LdQmomrb1uQTOMGfG/oXHvuQ49ocFoJ8/8Ix/lZQNCuCD+u/K78GD8eAvnhrPAcZh3Nu
vIa7u3wJmEEcWMU0ubZSgQT8m+2YL/0QUCtZGV0jGgIGxnyKpVQp1JUUlqrZ1rBHNsNyTBNUixoB
4AcxwnORubK0HP6IzKj8oM8rK6GVtNYx57CR76gjWohm2LImLw9O/xwQ6WYNHjBnRj1RjHQhOQJw
bIBSBqys37e/a6Mobf911msktVpEyBHmvll55vjtnM4b3VymGC/I4OZeeiWY2p0HZdDoWEn/oJlx
vBG3T8UviWbdWAQfkEYypHOqY/2GQDUgE6ZVtC7Fpia7ANLJGpEShsfSxpGfWyEU5aH/VWRpiKZv
90V9k+Y3foE58zEDuM+cXaBn4dabAPNXNuzQ/2+Tzk5YMyTN4tkdotI6zx9zellIP8XBKS0VzMwz
O2LB7xI5dMngECknB/rtQWz60wvp98QMz5E1hEwHvPE0/H8WAU04BzytHosBrUx7yB3jxO6tzPv3
QQ1hIH+3pLcIzOvyNcVatOae5rM351+7nnRy8BQ3YtUg6YVt6/t9KHywZVF3zQzHa42dwY8wnlYX
KUNxu8uhtarPcqrr6ZiltRi/wU92HAGzQVt61Gg+BT4xL4bAdvam5CPivnj753I+iZgsye5zwcxz
YZ5iWTmO/tU0F15Ma2XLZG7pU9L0e0f+H6EpfXA0imGoQPhvGwadYBUDRtMSlfXMUh03G6FJVyYM
0yEzj5BmFpSry0I9zx/UkcrFRzH58bj5Vx/z/ZmAsLItesvDUE0ctpN1CVf29VB2x3hrTfHjQZLg
WJ5U9vhhwM8NcBfQst7jO/zAiWfba3XOYLpJtBHX3zcqrqMocvKlI6cvPZbwyqQLUl2Q9YGTx/4e
/ws7auFfol9BoNgeuHN4iagFCiU6xTUPr4hQJbPJHroV4OA5WmL9/k7kGThkdFrow9TRwx7n03gi
H4eke1+mZ7/2HFUUlGdKqEjCPKfJK/nUyWfggB1sejPE+bugjm3FXwNEcL+JLq+oAzEzuknk6ihU
v4rYGpjX/oeEtijHRbPfsU9knBrPbmEwdH7jYBNXSQB1WwANe8mnswbL+C7OhoZKMxP/6ejxpY02
d7HOkpSyNKAqB1CZrAEo4/P0r0jvBbhU8Lxd7HMq04+MmCYmlu6ZTYmX5/HVaRh+Z8ZLbVViw2z0
0DUSVb1Uqxt2MSYVLn0oOXcQH4HlWhnrqjjzwflQWly2RWmoQBKe6limiFV5BjlE3QJiyIOrDDMf
3xqC/DPtqG7Qir+ySD9jdYuppuW5G0eBt169YxpX8Tjdr/AiXN0QDsStgeYA18+FOrITfNw74PG/
NTIoPeVNbTCvhMz9O3tYYrBk07p4oIWJnbAbb3sxv5deH+XBTzlNIn9KbS3mNtCgeaOmVLlVEutO
9CM4aFfCSP/6MJBHwymmkjWaqAOtk/FhVjXs/SdH4MtoYfHy8W4DIn+SuWkBW946DpDM3cJ6qwbG
RtLcWh8zHFPh3DQFTcK+pX2RGAjlymkhYRejJkhx9XazW2dFANAh+QGQkyPNH5d/6oeejsaQyuB2
kjlSWpX8atvDlsNRjOl8naQ3I5+CSIoup9QwGj/ZuesmDsg07KwtfHZ+Yz9GAJqUhUkr0OGxnBko
Wy6LBJSsswT8fJ+QSF/Q8z6U/7nf6uNqv2kQ+bLLqRWUtUkmoVTPASczvgfRXnUUuyWrmDQH7gEY
LyUslK8GTbNhAqF6uoK//KQ0v43rztYU9LUtF1jGe91TTHpE1+oaWLi+yxmONbaOG+6svEDiQxZt
Y/s/QGO6uuLY9HbJ2Z7KBBs8Z9wu1HBp3tqUU9PcaAH0k2C2Fek36ZWAzmJO2mpiBzraaYD9fx9d
wTY8QAfOSge+5p9OwMAuOw5QIMWbU0fMTdIHUucYhHb7+ed1djeyZNQEzN9ueRAuDr7NpyHVLOMQ
5qva4MTxX4Fc135XTdj+KSs4twA1sSdHg9reF++TpHYo6ChZhEGyqiRc24+lYTGeWrODFOL3Bn8v
vEsswAfMpSQZMlY8/CYOFvjPwPaA192Reeu7SPSdsV1j2+QthVfcGy4AbQAvvL9Mf8Z9+fXpFjgr
L6Lztdd72gnNtMCt4v66xH6nauY2UYMEyn/aDQx+rOY5OfSqDwZfzC3xf1taUCH3Zk40p/0nXjpF
ZBbg2VFTFSl58/wTf5a2Huol8VrvxpoBAA7Q5FvV3+gCYacxztwn6d8vB+N5zOC+pA9gEBhSEknd
hO/bmVQ5UDcfFoerLdJOVPE9/zXSwllgQGPh+cFLy0qCyq22lzEp0p9UOp5BJmcoKBTLfemUdqBv
dFu92P7ygLM04Jsl2dzMx46imXUhgOJuyjTt7XAeefvia6VvM7atOMr9TV8pHOkk/f9x51wTB7tz
lbC20nbouXgv8ooZR3XmXKz6ksFzvIK3YsqrVzMQCvQthrxShfuOMt5nQ9ylpxsFuGp6xvSQ1ROb
Zfpv0nARPYapFqEBW208piT/oPeYVslX9UTimRloSvYFQFYEQBQWYPYGqceGsjfVxthu/8DfekpB
ieWc52cgvpU8i7uJNkSxyPqFZGZ2qLgG23IfeTDcVVxxy9YsUkT/qaacsl3UNx3OKs33McSdkcsi
x+fUkAvWM5BHHMySLqGVLuHByOUhZMJA6S8jX62BRHErLtJfqzAULE5JioI2OMdJ07LbFTUPSZ1v
vNpMBMh4Z4XvOkZQ5BpRpsgQEsKMsat7KY/QPLc2lrd1UG7DuR9aeXMCel/ziwSHIB/0a7u73u1Z
uMEmVU6qAQDOOFp4az8jXjz7k3MqmD7iP8ht51hZ2VmQxSZtMXgrLzQmaWw2SuqvbZiiuCou3qOC
1pDRRzJCgXcNTD01jJrXvjLhDvPNy1UO62HLhFNuzarRGcDZwGOHzBEdnNv/gUTUeVqHXu6MyXPV
0aZx9NBGR0+xvXQ5gQ+LfBK3n96lXBqA6Ak1k4//fyCVop54fpzW3Aia8od86jDrLVWmPfPki4A1
GJrHl4WZj+AVqB2b6anrU2KuyICu+Rcm49lNARgKgdbBRUFfJWoHdU0OeloVe9+cBa6X/QaggbeJ
wy1v5ld5LX4/5MAVxaRXA4rxXUs9tE3WEVbGyDxaprSztaXs/3Mr8YucJBel5hJXSTiA2fw5n0ld
kwHh3zOVvL9vGFh7od6E2RX+AetaPPoSrcmUVEGnwDUoxLihEeMRYFqR7NFCbqFqNLyqIcduGnO/
BtgZBbAyWk4d3vKfrw35Vq09beiD1PhRhyxGJNzn27MARRGthksN/oENzOx9e5mW2MjcDsJzZnF6
O3lnIPqjBNOuACCIXsZDYUMm9C/RIXzxUJT1zy/QG/5aPZ0VFbifBPJsfDLLJr9ODWacqIKe/4hY
M3ngAI5ziwY77u3m/5DOt9aUlIgkBcZ37FMdW15e35uD/OXn0QTCkC9/lOOimpHo8wjXBgI1c8v4
7ZDHLyTTHZt6kbfvBZDPBToZsZk1Jt5I+s5WTScQiux6R3c2t97yAmQSFEta+m+tG3QSLroZqQ+k
i97NoiO25ah0JhlojW3eQFX4wpOh87EeHLLZaFhjMFKFiYjLvnVgLCo90bTnGDp9EnTq1Q6/SGXw
CkPt83jcDGYLTO1rGfDse3Eucq4c0EX/WoCWmgaJpGl/omc6vGyCXy8j/urnN3PW89r3ZIb/E7K1
kA+zkfSfCBU8I7mXC8lnBNjmSqs1JUoBV+o/9ZeZjTZMLh0aWo3aO4SC3q06xRTW5zfH7GgP6bkv
CYCFyCr0Qe7/FNXRG8WL8mazhuOqt2Y3tXPhgQKaw1nD9vEkUZgrR/tAJkVtqZP6BTX+jyFJIGlZ
xZqeSzUN/9ekSsrk4ou3NRcXqS8K6XO5hBQWwBgP/J7HNmp6FPLL5/EGp6OkQfvHEUm+NT8sswk8
LW8/NSWGxyOXC5/9k30kE0VIMfwmkYJkIkEsY8czhgoXkFfbt0Ec0Zf3js6fC+RXJPYgCcva+Cwe
JW5LGQiG4R5dUou21J0+BuHZwwrI1NHXlUse5WgAPY0q969vNy5sUU9S6aDCC2h6MPBLymvmR7c2
D9Mxpj2ckxBe2TZDEJT3NXQCg0b6Tko5tNK7DhlgHdBPljNHx/oslHcjJwPj2nbOVQiz1H7IeC+K
TaHkRHStg0mMfxjONDDNLRu440Vsqk3A5ZefPwnScQ7q7MxvhxetRJlhcai5YHWlwYU9dr2XCclR
VTpighmDg004fuUbdnxXeuemwCvkD86aYsamfUJ7dmii/uYi+TOIVIia8g7qygZVGSkYXAyl4lAz
CxZwzRqYSzZ40mdGUxfqkg0fOR5iKBeW7HtIMYopt5pX/Ppgv9QOIbCed1hM6YnB41D/5Cxv24r0
qXKyvWvB/k76W0kXGUdo+67uTrLVnBJjGA8aadeL//KQx18HIjw3fS3PiZ3Mat9BhjDPbigLGiS7
JLKq8MQYUW86DkNMLcpuYKY4+jWiQRTbTUoWOf6kTBbX440rK0FaTd+6qtlLksGja1oUmNXE9+bh
z5GkgRInrJZMLID3f+/teDFbcGsUz3X56fP3tRoTWNlIhqSRLauopcrFPWIcEjTtB77yHkMHashR
kQ75v/Pwbn/M2opJ7a2kiF/B6UWD39BI2k0jcT0OsqyqMkueqM2Vy1/CYkcQq6NOPhUr7bMaqYF1
LG71uEH1OFd7Wy6kOaGg9GBsaayk7xlXKP/Lueb8EI1po+kGmtquN3FVqyMB1/X4sH7ufdgyDuRI
nWPQRL0nfLqbjlbkz0tZoAP5h/sitpTezvLKng2p6QABLN9E3udLV75Y7/+zzxvWh+Dn6aa+DhCC
5io0VSoJACV00ZoSHAlLVmPTz4jJx/SYUwk5IoxsgphJhvd2gcLiqxp3I3vqunKuM3kGJA/LTR8B
OCjTyDb9pBgFgjGEOg0ssnPlBHpqY0NISBPKnJta28jolKqbC+raytfEnctsDgUDskauU76ZLWi9
UMwh/S0W2EcgzSZeihUc47HlCrJHoAUHOXxzz5ievKiKzLbwIBduSgqmH+xpUHwTl/Tx0rpvH6X6
fyWpWvmgJlS82Ct0F0KwT0lJI+TtaGEWonmYXyAaBzkAxNnYWP17bYSINrqJol8Pi1GXSVJr7MAA
JrlKD8+KjCoQXESHB1FOLuOFWUetY/kmvu6hS7ezGqR/K07FHOM6D/lV2WYkUzz6qXz0ZehZdfl3
ZjWqoeuBYDPH4eYbFYqSPplaUKtY8aKPFk+0t+kGyR+Sk1VrxQJvfepjjXInSbSE9QLF4bLdoifa
AZ50jxhZLt/fWs+j+INDpSFNTN5cIzKIDEHSYhKE8mbOjfCwODSLv+4RREC8uQ8SRN2hsORj8XCh
h41jJz1k3prVE6o6pfxAiluRcv8+OFZuQuxY80Qa9PXR0IkpI6fqPixJX6dlI7S/cxsDAxPIUByq
Z1+W5VtaS1+zhtK47lF3WkKh7014o0X492yzeg3pfO54X3REXl52y7a8XRtxJbVsNbg30VIU9Mqz
uA5CJHiLWOn/pGXMJL/JPn62Sdv5Rh2RZvnWvBXfBeW74gftKoo/zuEEj/sXHG68ERsWp9tjemwJ
KmV6cVacv4Hr5Qso+s/OEKOlMq3WMdK4QjwcXlmVJPuY5A3OJsqYncqMn/rwvqE6TfjowYDu3HEN
fEwmO99F3YDy5J67EolUHep/N+S9eV0zFpj3b+sr3bO3kDKJMuOLalk9XYBQqPQP5nBZQ22PGgq6
zlzKDkTmJqDhdlauyEcfRF+leWTrBiLJF0LzP44rtrp8E789lQS35po4LOIqBJMAKkkjHyRyCAgo
XNR2aeRKTupePGVt24a9qq5XmJ5v8Ej+uS93Zj4S3N4tyt8FfmM0N9/vqhvhMjCXkbP2/PH8CW/r
bOjPXJ/cb+XSSYiOs3HOfVC+GFUoMRL3kUtGlQEgEM4rESjxindjnNzG5ZYHZQbPFwgtFoxForUP
kZLqWPq6Rvb11ppmXPU97evNHEDBS4QnX/+B0uR9LrPjFSnMhzV0MsLTd7Pe64OGtA2TIgAxG8is
GI267rf728tUVK1DxAmTV3ASPTyCdU04avl4j3Lh+svmNTjEyWHY7tpkPKT8kYyNpHiDGzZr5uhc
xIZvaYS0Mf5SZeIi0ZvJC6I9x9Y+O1pcUKrSr4pMxZMNcDo9Yet4E3Jkc2/fdO9QtKHAuJfATxU3
PCU/YIRu5uCvQRdc5+WxOKQYBQhToB29xzp7QdzqPFxXqxFvMOi0Wr/myo9bZoYiIkwBVa87kToc
krzYqE+7iY7Wr8LWlfwgm3FghlO1kZLpnYk/O6LM2Di0VOBA/yE68OA/YTG7C3M/ZzoazmuU/i1d
f0wJqHr8d/tGdkMKm7tQpegF4WFSVuHFNLhxHDXoybHoiohG/l2LkPKlFpIS+4zUjHVSuZeAP4DA
PBmsQR9Nxi5JXS4HlzZlCWZmZKnwUA+4H4lw5bWDGxHPG8eokog0Rqj1lzObMEGuQWCk5cZ3Dad2
Or9rBumFoyx4oEBpJmpA2Kg+rgULeMu/vtjm8m43ogpBR9tHe5cQ3gkRMBlVjBQ8PFUOJFqVq+sn
vrK75ftRlHd97xzVLE5XRu+uBPsGpOANoC9k6GK7J1cGVnOgEEXcrkw/vljRCldLej/WkJke9jas
xbJnle9CuonHPdvQumUOe/suLqiMIdCMt2w7HA2JXSe1t60xVInNwN+fvLQVHbQKdT/FFGsEZYHA
CqViwcl8SXfVIRM5E9lBQQ1+BqLjrzDs3Y3FmVhhsiGbRru5n9OX4qj03hBLfBBR/Qd1XJoVvMSE
DJwq/QLTTqxIPfKpAA1s/TvrtKm7nSXTORDkEOCXr1AQ1yFGlGTifRhwW1B78oSCzg/7NXz3zrYY
uY/B7/sm9XchP861Vl2AVEC5SEgxrKnqT0n7yNn+rB1u55h8et8MCp58VwMe8IO/wOP7Ot/p6/NE
Tzq9B09puKCiEahQpoPPZYA7TqgDQ5DWGatxQGuTjDZd26ScpHSn2tJtgK1Typn8x/5ktNwWsH8W
3JSKFba60tFqOCjVwjZ4pcAqx9uPdl7c203vEmnNNjKvcC/pzvAmdqrIcjg5evU3UTGQnDZz85Tv
eX1VjADRnKzsWMnLluSpRH1uVke2qWtu+P8zopo+WD3/bLgJ0bJVOU0M2Vx+ktcUtzdCSGfBczDz
RblLldRqfxdnBckZm1QOJvM6zONtTAR0rPz9TYa2SQx8OPPlG1DGFyBZD9Jy0HOErHSn6tNm9VlT
WthvNEXFz2uyDDiJNuxyl1cmoQ9CeD2UA/lqhb15vYS2Ue5dbMqiGs5Lzhki3TzE01N7tH42uAnA
7JPnpfHDW5Y1HtSHwicdSMLeUzNG8chMzL+fYYP5SEQU3Tdp8Rf7yd9PEI2JcJRkdy2iilfTsVOG
hJzRZKTTLF4NOhq4kmjX6Gjzgjq4pf+QsrpmTHB2wWTohxMyn+dzXjHOM1mISxd/9KAXG5nwmiEE
BiVa31MyOfNOCTa55iPn5h/ViZQ6F2SeMW7G8HehuWEPMI4QnFW7OgQvHFOEoNvshKH6QnUMx7eq
YLfuEB8l0a0zNciWjDvDbuZyf7cXq5nJsCAruuwLM2E59ZSHKwy+5Kfux5IW9lD0cLOhyHxo5ORx
XtsmpjdR1gfJM8/5OAfmp+mMkJKdR2iQWrx2W7e0GpFcJ2c+LD13/EUHKZU/8RkgDCwx8MlRD9fI
A5I8RJlR2ipV00TAtljY76Rwwb1ABMbF5fiy8Bm9rr4zdW7rdxszzPUE8Oxfwek9cPV50tIQnu8F
55c4TZxHDEmc/w/the4SHUJbjM+UiUKXBZRmAM2xSn14Z0G0z4Tw8qPg4w/V5nacvhn8cuyx4iSG
4KzbJykoToobEdrUsA4QyTNBq14xbo6s1pVS2QUMCb+TehBTjyUqo1XPsscbiH67pK7DjbVUkcM1
zkWt6Vimh3D4I1erR7I8XwjjE5/S+OtIsANwI0mejvSwg5I0fUlJQw6ZzeJ22d8NyjfzARqPXyh0
dlHfTEp//Z7eXNvDHBBS6u4/fycCisN0F8e2Q4YHineQ66kiA8T9oK/f4UVPFDqx3tQxl+NJ692d
ruXvBklcAABt42A0Vusjz8VALRqDcWIKAL/LZ5L1ivipDbdXhtSkzrvizWjFskg9/J2n4eW4DuvG
cZxKGcaswqKCBeRxJEuSQ6Hcmj+NxVtQ3BVeL7L26ITutH2QcWV8jThnD2NVYVH7xgRssx11tKJy
ekc6LK8s2xQLGmbr89G4S9SlfgQXOBdXusPVbxyxJXvrQzlaYvBVKlbI2LeEr9eXjDAlCXEs15NI
ZYnAWU4se4RQWCTgn0V5teWKgf2zg2w4+Q9xZGdnSRw6zPajd0uJCja3v89Zv7xR7mO186Lki58r
fR36AxFZy2Nn30me7L9fI1hzj2cCcTubgttoCnslurSCnzmbpKqMNGVYfrT9qn+16I5fOfSYA8qI
S3gbywKYB0NxiE1n924wa8oNhdDWqyxA7lGNzH86zidbPkfHwFmlO/8Rvo9UuxT7oWpIqrPg03C+
2N4LlM2GuPip3E73zVRacxu+/KDuzP0t1YHoEgukColkvbSZrBBZE93ZkEEWg9PfOYqFPdeshXRr
qCF4nWJPqCs0efrTt86m4yPrunjGQRYtSZ8a5rUTqotKHLCS6kZL5SR61MnXa2kfLB7COt23qtkZ
fSd6tcjYGaJpPdHZI3boDkEZtP6YHKke+aMyRhb/qUlrHeXJTxGX5GYqSN48aXSx+S0ogRhbicUX
qp82DpuzIh/8eRJ9j48AXK5IYuYh6OLGPkquzzYibsm3C7mLiVn+ryRzCTHz0jfsTeyzg4kXCHL3
Tgp3+kJdM+RHQjlRrMuDkfV3MIYcReWYoj7WzUPQocdObEQYlhWZ9Wutcr8wiCaZ0nMA7miN1fHx
2F/oRElKaKpcp/A2Rfw4E3hXHJoi+4aPZkRl4ml50xlfZQpdFQgMg+xseQYcUrEbgiEzf3buUXMP
6Amldpd/WmBiGGs8g+Qsj6jurWZqtxLZRDLPTeBx6iDLcvi5rKV9qElJokKRaL/fsP6TGUbcpPDu
1WNxKIhAgvJPW5pYdWbWuOojOzahvO9swKMAyLlZ4dBQlwWR9GxoFf8ZBdaEuNqvF4DpVPz/vssx
LYoptYrADLt1PnsOq6KuoNYHC/qNo+cvHpaMt+tgvU7fSX8H4P7PnWAzFzrUy6C+hKLlvhWTdawi
xPxwi4p/BkspAhDTC9M91rO21q+EyU3siPNvbdCwURnaBynRhft7b00x+FFDoUuFkSwkhb2ZOnEV
XVZCRw/NXHi5rdOFBQHv3NnMektMFoWzqGD/wOlfUe12jUx26AYj+9vX7O0GPw+O6pm1cncgC5jB
6mOR5xalowN5IhsrjvJqLrUA3sniRwaiJ7TaahFmAwuo4BgRyLjK6OYYToo0hv3YXKqKbWNHqIxe
SDa1bZbltSizK91dq1Arazx8+VGspNbVmKjeF/OTnmCR9164s7Hp/JDzsC/pmWM8XrsFZ2cHdDLo
6EHGP0DDq3ny0qT0CDshBPm+AMDFZqeLqNFPn2jlPoVsKmWHs5LFa36r5hZ+J08qMbImdLg7Shvz
pgPTG8adQ5nTYqHfDMtUzC/E2k2f7hm62MUl5/Z+7Ns349G0dkRf7vjaBFGamI7x2kt77HkfnyxB
/DlTFfhEvxmPpHfk+pZ2zL8nK0n7zKg6F8RISpbvx4g0QruyZZnVUKtLAvZwAuKn2LMTxQSFlpYe
JGcBtFBBXmGCZ0S8NCQk2Nqtque84zLwxGlmhvMCOQe2VTzAMMVaVfOswHs5ece/EbHdew7SjzmG
SUNOmc4MqY/1O+s1t2uQnAOc6e0IlydnOhPvVlq5UEx4aV1EtNXHe7+oLE0P2ipQvh8aPML3Bn16
LssWtgm4DEHdFqaf4SJz4rgOYZx1hQ6dn91e9RmafTSZp4Cd9mjZjjKGPnoauUXrzE05H2Vgrx5G
A6uUum5NCNVgMoSNZFDAkUsrJW4OiNrMqRDdjwTO4UhpkzjHeT+MwOUOTbTuqK0pdwbIgliz56u6
gca12STNSbgzBY2LLM5fmxurI2SoaogDj9kAgom+Tfudu9MMc2SHGGgp3rZkJ77wnVA/RUj4Qj1o
iv2ZHcjbgEcWqsKyrsQE4KzP2xStwXPWeo7WsGmf7K9n2t6E1nHDiWKUo1ZycBZWJVdOTOBv65/D
txlHSWzPxbx0Afx5RgiMZIwNYh6RjmsMFaQPRtWn9rHPUbtuj82+zsVOCI1vOYI8rS0WneBLFlX/
FMxGhy7WqygtME6bZj42ARAfApZphGGCMCeZS2hTg+y1tvMx42rNcYU9GN6QI3ON0YfpOCclNpo+
FVXEezGjF7z/ItkaFnK2/Blm8UfrVsCyTVcRoNtEbnnZY7csuc+96Cl+3OUmqI03rkr7SbBDI3tc
D77CGr+6iKl0wInCLhqv+VonSV8REtQqcrFF2yWAp3NbLP5w5rXOgkGtKytKTclerPU9us0pV65R
8SSciuLabLSyvZDIq7I3sZ5SNaR3/3v6E8PJBV6LyqjBe3Lx4/Pr4WfhFssHMpPRp+4Rpu9eAXAu
vGcNAgdWisbHd+ieTKY8Aq9ygUjvfEWO1t3c2R3XW5VnOaXpBGSoL1izPbXsxBopy5+zK+HicxV+
dNjpBuRaWfYVK8Xbuh8Fjo1516YHKwCyRvET6yNq73s4qxCBN5TapqUn4IBu1kUtnyVAuLm3lBPW
4U7U5cbejAmXnPSDP1CCmJ+IFB+8mdtClfXfTt69bcYh4mwPCJDZzFDRoMHNBDpYcw+RM22rRxcn
6QsNqti0XFUBtjjfl4hjVVUoc6B3tVWm0k29fXswmy8lqKAqt2EpCafcOEJdPgUh4BN7nKy8/xNT
YaXF8DbKMOjhjToARfB0c4x2YwxSPgLK0GUhCoAE9+xNxIsi8vUeU6jSg40NZ09Vdeh/uiBM7PdE
++bKsXtKnBu4/+8fI8TDYjhQbs0HlmTugw9ck2L1HO5En244I465+Z/HVhBruQkKSgDfzgCDO1NF
MbLnNM3pm+zNZpeg+ua2Cbk3cYB3TTPn4o9uDiTLXBW8j9qKNFwS6ypsYkywvqQDpYtG4Jpr+Vt5
s0/5asXzCSpH91UpR/0WFxD818cpItE4mbm7EFKMHBbX3jf9js4nQV8soHO4RVR/tO+2EmJjF82F
Mb/ZK7M/+aSSBtYLkevtvDfsbVDpsi5je4d3cylmw4okVhdoPGLYNa+KyKGkQurwRnNyvYs6ZYzo
pYEH8B/U+OYxLg8y3RdhicDp1SQXTV/t+0PcOfHUI6VayxZVAmH62gaS2Vhu60N+scnZ7L0wKN/B
L4qzRPv4mCC3Q4Z4jUBddbWd2f3uKVAvpewiqSbaHfGe9HAM3cQWtVrYzQ+nPmLw30kVyXZV0XSM
d1VcfGGxrTiu3D8HDel98RfqHeB+L2lJCSzqj9URN6T+WxIpjyqrRiGNxYadmb60JCV/XgUMONkK
7SwTvr4gOfHzzzdohaKAa+nUvfTqDhleOa3/btMdTYtBB66ed54AYFG/v6f9in7fQzNH4USb4Aed
2yq+4BXroI9r1mzegaWSv41O8hsjHwmbC/T8C8nh0vbC6HWVb3ZJM/Zo5pEKMXa2lNpN6QK5P4Ua
SonOiFo3ZydRDGoWRpqqKJuA1P9hsa/oRt5bQRLwQ4BruIEddhCEejXSpBnR/ybmp/vexU9kjh7I
vX6nLaKlP8FrJ37aOG/o2PMgAxEiPfbx9BepkL1qVSiDRvO0T1ELKSvke5MQsjSVZtXl77O94w2g
flAyPyeaYEBTPodGhs0ogqnzJ/MsnT/DqeK8LzRUhv9vLuuB8n7z9pgjCQJVoNgw+V7DTaYxwn1t
wcmLr6usE1T4FuXS6Nii5Kgz/FOTvT+fPgnKb9Nf4KSztmMwBpVSPv+p1jGAmGuz8maxXOfYgIcv
HbK3ySfJzui/FvZ8HwZX1j9qKjFsqJAMpHOGl1wRXclUYwL9sJiteUr2YZAWGzM7B2DmEN31zVKP
i9ToANIa/byL6wegtqDXgGlYkTZD7Q7tYMOsphcFP9sDrDB3GI2YX+jjtBXHaA2nH8BRFsZ09d/P
f0H+lsqw5FrDJJIU3u0ZFp7UItTS51WgONLQsv+w+Hqk77p0t6eAcvn3JKUB5o6fNYuJVnA24cnp
YTC004gEvOJQIRPpi6kWv9zBoDJNJNaAwkjDZwjtgoNjEZmKog2WRIVuE4zRX0GjDnBMmSzUy1lu
h9VB+C/zaRJMglg/CVtotdZNCgX/3920FbKjH/7hp0B0TjGkdiyd/BCoP8bko8RcEn5QSokP5qvh
25DwAShHvQgUzFOno8fwOHfy6wZTvg4iblo/jRgadCGXtnmTVA1kcGPdchGJXkNgwEF/dnGsB79q
HzZxk6EfF3RIcoQF66geCxVUwp6yrp9WmkBm3RXxLkPKV5mwKbEYXd31ozuvQgeXPpRQKdMcSuYj
hiymbgk0v5bJkvqfaUNBtEJ/XgN+I9CRcxmCxhmauPhHb0fius31MjYW4Igebika8ZssfMn2l+l+
wibn3tZhAxCD26ZEqGJ25Z3QPya68RlTxBruhAh3SAZgOGwPQ0HqPkTiQN5oR4QFoppp5imWjzeJ
wRvGe+xsGOANbB3/yLetJZz5/zHiBDGylkz2UeId6clD2gNOVVHp5++sD9sCDCQzFW6hXr+B7yu+
wmEwutVZR6ueKnIscQgMTzTKlGdhLwG19/0X5VZf5dOlEo6KeqKB2Oh1W7q95VCMeQncqdOgwxj1
a3nt3Xsb9lbZ0RdLh747oHgmjs8fNqT3Ojh3goVm9T0IReiE7FnMEWW54HuLt87m0isZIKevau0S
798hbwhgRllZJEd2ucNpJT8Wj4R15aV8VBSvkllVzq50EX5MyobvfEwKjOI3pGt5SoduLdYlroM0
PSfTZBBRUnoD4YUEjr+Apdb4BWtTVys6u12u6Ze9fpEPx0MYbwh6p8nAmiJxJPaXv9UdeK0Oxl8I
F2jhiDtZOqiqLO15nFuoaVgntTG1PQkxsDW5WYSlpiD3OeZTYiewnhLsOeZesjNMY0IqfsuwqV4d
oqhsESxrFrse9YYHyGdn2z568Hv+ojVxS9OSQK8kJL52P00j0lusidnPGT3slOr4QHrU+PdlNlXk
/+mX3DE0wei8HH0RqTcMBy0V1grZrKKhAdBeVA4kbXJe1bwia8pVZmL01lVIU24c6qrnthzEmPjd
qYoXzi+Aw39YkGS9H35afsJmyFRzSp/mpjCuguqHCkiyvSr5flG4MfetNU4ZSqdINOR/w9UJxaRz
jigSMqWDOXrV82yC+8TzM53/6V3GP68aN0B4acKzlzLkQP4HlmQx0YNorIyIWhsYEiP2ub125BSp
1OA9r6oQMhF4oZaZWdJ4TQoDy3IXui3vt5wmpkq2Y+YbATKkIrjEd3hieGcIzTf5BH7tempYhj3z
kc1s3n1y+6lLfo21O0s801jQ653pkpndo6kwGN1wtE0WBO+bR1HQimgV7lir+TSVmXtVmYJKcG/C
2NcsWc8WittDWFq9ZankLH4+SJvRDgee9BbcbM1PR5p6gYg/W47VpuhXLpYxzh5KWcDfZGvzztCc
MEEcudHAEUEoqvR+RtyUyaYcz9/FS9AaI14+q6ntAIhVgZQ6WuEJZoEDe+KJVCAfiX7lxYCXULOr
s9yxL4dA/XNYotu5R9O5mTXG3SF9rKFf8gYSxhf3IdvH5tcN2erqs1Jo2ip+z/TIBDVk/DCOcSm2
49vbMMlMI9vwTW1BLhrhy6wfGK+H3gwSQYuEWWknYnzkLjUm10JMKqF0vriM2ahW7LI0ju61tZul
9v+VEBclh+rySNFNDJA0g+tDVmq1WxXoTfFQL/etJSed4uzEW++42WEi24Zw4g2OdJRwQVY+J0fl
VhuQrb5ruzEwg21wJooV3UhQl0RabN+tYDqBLs7UL5BgTxKXRgq7S7maUfOuvpKmCrDLjg0FpuGq
QFkq8CGV8j+i0wVlN/mJlc7WRwA7aULttz0QWa25S3r6AJARERiqay3LpgY+kCIUG5EiuQRGFDJw
tQF57FFkKSWJD1HziIxMlxp8Cpxk4Q+n9tMKauO9KcvOs6AVddlstvgIEoFEuUuIr4a3eOntYLQF
/+0G9eRkxTh1bY5XSmu4ZbdACQXZPepIdrjQkqtzGN2VMjI6ZRcRmegtrmOUtDW80WArv942shde
see9KBjLz0Rl9JpFNVDbnKhKCSYNgVC9H2JcYgI1yjDYekvgsTT/rnHzmtYCTbLadn/VZaJ2ULU6
ZeRiG/1mRsfm6EgBtjYHDxkkJ1CjgbBjQKfPV+u186Yk0W+Fk6lfVEU2I/KfiK0zVtHylnQqCfXu
7tzHjhSP89GPvQpy3Uj7bLb9428jDFz1ilGWo8SPUWJt5vPDGVT17wXUgSgztPV2jxkf6sDQI5RX
/53kgASemsXH5DVfoFzX7nt7mXfKnQF7VLCrT4lECTPingwBOjBvL9zNqtnoYaAupsX8YdejEpNc
AssQ4LLRDyw8gMeHbkZMQh6Tl3D3LkpnkAFeS5/UBn0DKPjCi2GHHWBlFVsgNPWQ9ShUG0Od5mG6
nZkw9d6MbgyH2XKevwIXY7E0ag9G9suY2kc6BnYfljqpKJNOZe/j24yVOlhZm4Q/Hk2IMx/TMA1F
hyHzS64arwtyV8jIoFRf5DdIvchUCMxmHirTo5xOQYKTcSGKgXIYByuKxlJgUlN+Sy+nC3IUfDWH
V2gbsk5Ng6v8w4qE/wZ2z1pEuux0HT3OXixSew7MF+cdjFKEG/kUkeWJsN8k5lmpJOPqSkexUDLi
iau3syKd0L0A4i2lZzqwDyGmLu/zM+bnhaqSf8pLBJu40cUM+p509rguwvfCtu/XKRCney/y4kJs
Rr3qhvfWcKOjYoN0yNWQRlbswmxWoCVx12D1NKpCWBmvZmDI/2yS9QRMiwERcJIS4IofkGs5qwLS
yjHAsn1ulEh5SnKV3o2wYAql1g/zL2TMCAmSsyZ5agG5hUJMYV+D6cqJKMRXHNiAu/scYynO2s7C
DKvJq+iucF3Fcgf7UXY0nGPjwtU1y8H66r3vCk1+Ykr3fZruLvnEGbG2IgLQWMJGqAmjUrvD2xmH
tgCf96lImC5uz23ae+Xp4lZo00+j4c2S6cdjSk7IDTwKykOcMC14+p5rmRwjS2gDYpiZjLmmSQrZ
CcURfu/Q9WjqAIunY3b90xAn+xp6SSsH+MXZa3YFaWkMLgHeVFjzw9wzF+hAQB1PgarvZFb0fwqp
yS4lVlGZ77chkarVi3F1i69F9V2xiF/EqBqg8/zE/h0H+q77uuAwfNZQOI4BjQNx2QQrqrNajMn7
NmwDz3Rn8BbNzrXiYm9v0d0lU26e7rVZJq9n8MiYq4O4QC6mGYTHmsNgXM8xBrnzYfN8gFdqA/UA
EnQKlbRlnM3W9EwzVyuhMUMQodtrXfXVeQ+lLj/b2YgqEtrIiMgwGe3S+R7r1m9xrKOUEzzIuN/A
WJ7Uaxak0YMVklc3I3pKZBUPQJqEEY7FCOwGr2hUS6Tr+sB1AG7JU+uXimIo9cyVn5xyQ8hECG/V
eefMRyhiRZ4TQYksx2sEJMsZ+ZNC9MkZEgwtfO04j+VkvxbjY4mleM8L/uQ5qINw9SqLGs8YxeLa
yO/EIE+dwJfxPGE9UYPlgH+8h46I+lIqLskLc0wUGO+RZ+w4hu82NqmYHNA5+UWjq4VK2p7uDnt4
myYRP/1xG1hd22MxX2SPwZD57r7OIh5TKLjPUYSmvsgNYK0hTax+0xFW/Fr9makuG5SYVlFqbD9h
Dz29KIKuzXZq6hOGYyFuQTWgkmOWz3krz54BrD3lOyblGyxo8+NFusqKx9rZuWVLsBBN9u3vxsB2
pTAApejn8q/ftbwJzQOYi79kxLeDiksV6eLaAnu1TDvwVkigAr0K+Rk5JvOYN5K6ALWVS5HaCt7P
Q13xQbn9lx5LVRPN2GZ2Wylj7tmAhFxCNDeh1ykWExjmR8RragksLB4rM/tIqZHqBIYs3Z3VNuLL
saKjnQ/r71tL8rZrGb7rBIvrOWO7guY+fq3IUV4bgvSg9N4rvwEwVOxPKMK56d7yhdygAEkfdmOG
nmNYzEqVT3sRP9ToAug/c34oW4exb7FVYp+9Qz0/wBgvrKrmwqPNp0t6hKf8og3Q5t33vb34cnnv
YuFUDUX+AxTid8CWF6BGLWzTWYZwAO5nowb873Iujh+iSoDT8ucVYQmnQj1bKXhecNPSGDH6jbVZ
qdSs0a4dZYPyTQO7vnlycMKYghHaZ1eiUDsBVgTsnzPKBcGRAJpyE8KyOSItPhHkGXVHMxTvdM2f
p3D5WmTYtW48pZBCTSBwf142Dz4Exka/bYhP5V/0ClPv5FIKAN8PKfHWHtXi057VzPbEx7645yp/
xvZrWBF1FtVL9RMHPN2B3xiWyauEOkXWMN6gUT4eaR7B5EE44lwSlskxeu2dWmYggnAhqGwvlCSE
d2IEPNe8SIKF5dyGkrr/ejKD59F/9KRsBncW95NldYbFwq9KbCyP6LUwz7hofykohmustVFKSP8p
MuyMtQ5QxVBJFJq70tQxSaNEwW22o2n+0iL+umNW4uvcAnLJ/FWBiiHYoe+Y4wnPBw1hEcfWP0Pj
zIQ4N5SrvHmwVStSjChwj3dOCbSkxkgyRxiDqm2pmaa8CKVvXlGVOBjMfIk2xzubeiaxcv761x42
tdNuhOTJfY+LB64iNBJd/QqSqp14GaxzUeWRQqlorKEWNo+TDk/7oBq4IOdzSdQf/6YWxBjOT4lq
Mi5QUxn8DQXLNYgSU6NIX/clcNpiQnuLUDN5jxUZr55BUPsFFIK73FeD9s9fuDMG3m0L9I7P33GI
o8qayl6pln/eH9kygV6yKiR8W3Fb1vV23+gWnmTbGZZ57O+c4Gu3AK3FPnd4pC33PDe7BXl44oJr
hn5GfEVINYt23SEad4GM0/adikPB5EMpxz+MhqrBwqbcQSLJHE1q+xjL+u/xUzL4ELcpVi2Vp+ua
tnyuea5O3AN52hBdQ+smdT0kfMwin4Y622uIOoNf55IX8KH+BW8fSUh7IbfWMh2l+p+h46K3lpJg
gLoepypwnQfltCqhf/FgcOSo0Ju0czZlmZ7EfN6G0lYkmKduxgHgeCDCXeaAQ34u79iLLCJIHnjh
oWuYSll4cMLeyjkyhGgbqTsxJFFAfO8M0ClWavjKU4Vy6UG7JxabTRymBZxkEyxYkeuA4JQPvbei
WBVGxggwEds16M+dFgTeXzoh4+IbsyVF1BuZzi6H3NPzYV7/HwK/XXcP3Z+292uU1IVlOZXsze6U
w4PENYRPjusEirBB1ewdOqR2mkLQqHk+UOajd034iRiD+v0qzx4xt3jLX8iMFdFaXEy4Sb13aXqT
DSat7Fhr3ofqigZH6RbgDEZ+nwBrB3KRZ5zTyyBk/NIo9R2wFS8MtHFq/LVv4eegmng0/Z3eQVtS
C87sDPtp4gQwurcR243iK6wSvDI4N3tXDuXbtpJteppeFe+UyMu7/N/RkvN6pZ3AhfnFwQwfBCvz
LsUAZzPWv67ygRpAeO3zxZtp2aPETZ7yMgdebY8mPIsqT1UNbpjVJxekHfBxznPYmAVsHFIIetsr
Yt5PoixmG4Elqqy4zKtGDZPJxwKjkFiMXthYhuOc+BX51s4mvWdQXmAYtsSHyr83NnGc6qv85gkc
+87Z2f/zxRWZ5jPo1GXqsPcmdQPO1PVAKDRYcguTKu8+DQfInEEoV1q3hYo6QtAecoFn77s9O6Fz
8fgVs2mP4Wls/BUFR//SUCLLNUUJbs+rVPoAifLGZeC0Cv8ecEY86dGGuAZX9q1vjzeofF7SiVVN
s1coJy/b1NKkr8iNdH7EHqAwTQ/nS2xW50Edd3sLcdiCjU1VdeGj1CZSZ/SboixOsw+RHjF7z8XN
fQw2qS4UAt+jqViGaAQAN8brMXh/mTqrA/bfdZeg7iEuon1gUco7ikT8gHT/VYu6NVWFfEKe/vtV
n+y5yDjwdu9feVXGy0+MlLoASTbiUifRmfL89iSo+f5KHcbNTaa6VIruamp9bs+gGIj5tZ8vQlRN
AanPIdcGQOYys3eDE3KYNxR5Aoq9pjN4+UReLBOjUldHzazFa66RLbLzQYAQrr3M2+YPE3yDwO1y
K6jA5mKgW/nY9qKjroxT7BV9LrpBwp25qMvzF6o46MCC0Pve/bbqfeew2X8QMJewKXlZrnYS9cFF
wpLcFKaxOHk6jaMk8i6cTDT5UuUMgL4jgrZPPnFOEXYTDM03XwB/NFFMaRweG3ktUO88mosIXPxB
awoGi2BX0ExsdNtaWFl6MHMGlaM/spo7cWWXHlyS8mdJ1PL9RGfvIQsh0PxXeFOHCKmLxeFkc7fO
m1AVRHofCsZQjDgnm7JAGYWTfYqOvnfxnY4eD1S17g2quShyfB3yVmj0rO+xDWlonanw2bfjuz3H
gHK8omX6/SNG6PDN54ZMTkXiu5Ohp4tflHonRC+NdkfnyLxQI9jEzOX/dyssoT2+/4ONskmlSTAO
rrfF0bbkKHDN2dKCYZI4fMMUlXyohBUahj0SmnSmnYHZq7aXVTvCES+i1p46d9+Dgc5AMw4UWikH
WdrmbXB/r3OVUebNwr7WYMPlInueP2cbt1/ITLPDZAyX1nrU+c8HUXJ1qX9Ewvyt4eOWstsqrkKK
6fvH4uhWJblk1hU7GJxKclFZqbaUraf1WCqsoAJVbtXoJTdrA4FnO0g/+BBq1C4rwqocJbFCsKcl
+hYahli+JCjHpVqUW++datfb0HFo2yFH6H9pFMOrGPoIQQdyhiVlAnX2zbr2JmdPcdBApYABL+7o
G5/3drDo3bQIU16hY2x2k8yd/izIQsCp1bX64o+yzbwREasO4CaRi3M+up9YS1EzHt3sOlnoPC1p
DoG/IBaSoLsWxYdHNvNbAwRjC7C45wwrFjKZvFnNGHd1vo1Xco9Uo9vpgXSupHASfkTzyKLEXBfq
JNfRW7DPC/Zl3gw86orwHLvAm8qf+Miqm/V4uIl0DT6njIm4FgtXh0qzLovcPcE36NMUv0KtKJ8K
nm6LXYQXwhInIO6j+gAgD1cOzEHSAyCPA1QAtQJVNHMFUkG4d8qtQWem2xWrVXkNOIw/xwzprmJa
w9eK7MW55Fj+nBzCP7iJoULoNzUQtYD731ApucqR7cGA84vhSOZ1xTZYZji/Y1JXa2EUMzMWWYr4
t9cKey7o7jsg+U2TL6djZZoBCCHY6kIbOr7lCxwV5htc7ZTdIh4T6E6KHBIGcfKNmaD0GAmFR/kE
V4sB/xPkAqXbLwbZPy4FnM5aJzfNYEvj6gS3zI1rsa3JE0Nev00YTwRxsbwchX7f7YGskRPsG7iD
41pZ4iU4PBBgA0N5fgG0LC9CYaMOvx1mWTuSCAEN0v2p69NdrAm+o2qbKqun8Go1rdYasfQCVUin
OP+TynVvuS6d/bltVaPPb1TtLdfI8ExA4SeInn2ceeSH3rwfHq64H2S3bDCD67rCEf5Ips7b59Ki
wtgoQAk4NJ6GOhpD0tSdJf/BYxVS3eB9pd6mxbchHsucMBRHYdKN7vuafNgpiY2+C2URba7BFqYo
OPjUIHy8SF4xsvQSkIL+785qwdVSY9XADMuJgXlZZYEB4mXOWQQI5RnHXR9yCtqu+WH7K6TDalim
XP40Mysva0D6ihfelQ/WIW1jVjGlar91LqUr7BbUrAdegAUH06kQGZDMb4IJF8yuQgaAmCDBavwQ
3G0m1DB/lFXQWkGIx6LsXLYho1zf3P03U8JyVxkd40opOA7UrsHtamlbPqVj87ENyid0zNb78geh
fr8QEXTY/MGa1PxvoJkKSH2NiLIC4Fy61uXM6/FVKKN33d/ju7YPd0L+/oUYHbElsIIDcsA5Fi2c
jnSGJ9aGetiio3HB96gAiHbi57/XR2ioUIgx+gPQOlL8FUMa2rzNpniCuNRH7E0t30CA7JdwNJSU
KgigxjQzNMStJl+uV2eDpNB9Q12UVv0AdsES9eFX9L4JIZfleEqBvDSFeMl9Ggt23OSkg3I95/4E
lvzzE5CpJLf+RBAmy/nZNhFuNyKM4I84IeHWanoKexpMngZjEBmXNDrcaKQE3hb1RorE9Zq26pWX
11vy6aR+RTOOQdvzXoarC4YJMYPdzHNXQpzdKHZaz2ysbKstoqBE/pDD6AoaJoJ5n9wfEnzDcqPT
AItCR4GD0hxS7KhoV2YLCXEwS5n2bDiiA6JfS+b3JgQhBndqXbCCRfX3q0k0SphkQvp6zVi/HCE5
xBjEUIg+WySwTlZOhFLkjN2mAkXtXKDegp/h/xc1+B95gUztLryMDlhrsiBIZ41nK+dNqV0bI54C
0/93eNaSt777qo68YHETYcL2VHw41jQZfI3g04aOj188unqYOxKtjOZ6AEhXNrv16k8qw5Mx1qNH
L8hUp7MEmNUe9ecI9dNPkVc2kUJyDc9CzZ4JL8JlK9jjbvSUdan7jw7e7Cvz4kirE/KL/yskCsib
AQw6pdlErBfPOpXwePx//XpCW0w1IB6dACXfasuDUlegiMSHIYnngBK/AEHmacsrvDXeBOnclJxn
i3+Zn6EmHUfWqShFKwTabCCaSoufFYg8Wz5cCGnsvf7aTlvDhy4p9m2evzjLrrqVBaZAj7iqigzN
4HVgz257Wk22CtjN71OWycgTF7QJqLGbwN1A+Toj4g2IbXPwNuKdOT7nweuu5e8aqKW9eM028LY2
Znst2ukncVeCFWTVuw+dPi0mcN+zyiFPMghShV9V+ki4hHBXvoHSgX1ylMhIwdQAfyJ83JSi9BS4
TNolW8p1G/VtGoqox2hAd0uaBTDAyghzqPF6MY8mReLPMJQi21ashx1S6CX6L5EShRSTmCbugeXv
hOoYpN+B8N6SGaRGb0slwY7M42rvlhEg3AXXSb5jiXKMLFQ146vImDGkqo5MgHZh1jJiu+N6YUe/
oLxGBpwu3Cd2FKNUMENh/yA9hBQGH50zKYiArPH2UNBEF4o7WsLJn25fgtArUytyp8pRA9xrWLDO
wSiTJhLY/e/60jXAeK8STacY3eKgvz0TcM2JyFeVZAhDt2mOu+NDoFxWiBFbIV8R75ZnIZeUP1Sg
xfufkZmoxLqMNYCBFCoehx66oKsfXvcla8U0puUP4w/DfR1ezuks+fmt+jTLfVGkuW7zsVqf9E0Z
/eRFPZsvVFJojHSvNpBsnZwhUUzpG37Bjf1tRbAlgJqFxvXIDQjYZ9MjqZ1p+jPoONLpEVPCkrhm
dVzdn+5FOKFTiYqRhC5oMIJFrpNeFdmQge7Z75WZHpfvNanWDj5Hsm/ZO3twz9CkO/bhCuuCuJ4s
kTs39uOPFZJfhu+LIZvIN3uePZAMnKSY7kxs8ReZH+aURkByNvfdyJeGmedrqMwrxengG7UDpi85
uF2sL8JpXX+w0s9yoLYN2KdkTxZfMEaAwNgoD2SOLmWzgTe3iuRik9RAVZ6xwmUWof6tLVHUGvSN
N40rUTubZuW3SikCR8dbXsPBxxOnXhH1JyRfmClPFEBsjvDghB++w0IfVkYfgF7cxtZ6gLRDKfYr
bmgze93izu4tyJeYVZAQ57zgYwB3c/bvuJsZv1VTuq7FUQsFaGokvctl4y3OKe8cVr/sWzpCb2qp
+pHrGtkB3JyElGZJjnclrrbtr/k/B9XOiSuzSdWYj2WWJKbxxh0yTM+worTqCxXF8SG1RXx1ieOn
fageG/P5tgwY4in6wPpLevXzv6egryh26JQ4eZseYdsotl2TD+gcGTFO1Ix3t9iJD/8GXqDVX3yc
WnmWb+ubGfg+Wmvdc2elZDLOxwQlutv9Vs+kuZUv/S2I9F5RsHrcki2sKf6xAgSNfUYHloufdsY6
61zFt85SqDqj0r7JNUSuToid3PL/Zws+viNqEn5Y9rb9ZOnq9vG+sAJdhKcr7deH0ndARPEijoqh
hX2BYOKmpAtn+vW3NbYr3LniQ1AXV36fen5OzWNoAFE3d/aQz11kGlVEhMvdh9AOugFnqTRmmqSG
MK5xroAdKrosYUBVEANqME3N7tJoktVaIK89h5PU00liB3VvM8Uj8H6ng8NAzz/yc5znBX9CO+Gs
gbxgfDozvOU4xci+qdFsEGiL289jIsH+WIV+wKtmF/znDyGM2szgg9RSid0giKyz6vpi05rnX3cl
ynv27V/vJ3dbV6tl2iKNr2AVsJsX8EAMClvMH6+UpepZkanIByQ5lPKHSFjl8Pi7KJOQwySrFPpB
TVkg0POwTX+H9JdLADL4hq2di0/YM3zhEAeIC+1sj7Y0R/sNuBd7HZ2htbHDttTLX1bgtUVgIljW
QsgjbmH/m7Nvz9/aUyBj12DKHkH8WrSZdU1Zp5mTsOluZ1yT320akB0kDAww7m7CHYcAA28ymGFL
kM1wgd0UImdt0X6TSGCTcj/olVySvT7faJpyRkvNlOo0GmNx6sb4qqq+9FHM758Q2YlDc7+6j7AW
kOuMvZiYURKjD9LX8bfFuPZJFfLZ/uVLFjscawUs/3Cg5f2badzF7khZKgO+/N33ZfttPH955rbl
2uoZDWWH/3v/zKAUufFZn29nNjo0FSKOZV5qxK1cVrWb3lH9nkbEml/nQC+1jUCnctRWXlAmJ9D2
AFqXFT7Umb8hmheIXF+8Z3Rjw4QE6W/4rJJFmwGx140b6DIo1Gbq+JiFKd+ECburiQ30joKZdbpM
78m88iuljfTLa5FJFCAFV8s+D0W2EnyueDEn3otwvULb62ScIbuYZAnaSnDtRbfaIUbGqXtTGBhb
g1Ho0hKNvdfLdB0Cve01xNTMmLb/FdaG45cc8ATmbuj3bPL/pBXFm6LzgFZSwD8riIfc4cR4kB+y
Sd/G96twjo+FRvu3yZq4EDuR1jW6TEZJQ6/hr4/aiXh1Ty6aTJx/3Bu9eHsHNgV5yyy4bHPzCnaL
78nxHj7u81pyC162jD5IB9HhYpQNM7cLBipSY/UEWfdT4zf6u5yBbx6Gt5Gnfh0S2BLOXrolgoN2
PVh/sx8GBgk2D2I6q+36ekO49lsSVo3bgiFMEBkXek0ctS0OrgrmjV/VoLU3eVDZwtlKmPN2nctx
aQL2OIDTZ2hBovsgNcR29MWiJjfAN7xcc8Vtx1GnvKsyIyvq4MB4OI+7Fse0Gj4VkwusO2oHJhhA
w/kcP1/E0D49wWMDYtq/fEMQlL0nTK5wYTmGBEDwGlm9MvSu5RzWfoU9CYDy5MEs8CdTAR7cyAd5
xJ31WrPB7lCk2QHDYnRtPWhMrGKyyim57ZpMbqcf/kllk0M4D+iU/GHTrbOLULGUve93G30pgoak
U8ErDA9qnaRzHQ9eUX9ie8jXqC9nhupwL8zW8DzAII9xDZ+8l/Hgquf8Vpfeg7K/IU9kr+ff9uPa
weKLGPhEHgIfEma9W+/nB5CJV0xpk6mrIJfUusZc+YHL8quICPfdozrUSD+OUc9shgbFgP6W4WCA
4mR0tIATdrExJb4tHoskjRzEd8mfENxlZ/i7M9cd4xrMRiqdO/iL12wWoi22oIRge2zv41ykV6bj
6tQYkCSJDpncdw/WTeOENrTRYHJ607cnHWVDK4wvMUnbDtnaYiX15t2uRkDCGUZPBqEgfsXX/tGE
ECpy05T/Cnf/P0TzKOqfDU2wHUIEFf+CJ+WA0KcNOHvC+3s96aM1X0/6IcPTZtqnxSJLT/2Ig7cm
iaZyRowG3N/dUM2J+pPyhDDL0g8ry6thcWDiFoRFm+v3ZnZ/QjZUgCQzBgBpFqTV1O6n+x/Rf7OX
iUBoPEx9sc3GJ9atAlXOubtxV3oxCUH3EKhdL5/cAwSSzK0Kpx4fLQlsqjiGoG/Xdz9YaCAVa+A6
EaWAL6fzl9+veI57uOMIz51KLWd/K0JVoJId2d9S4yJCTlz7gkDkOdQjqoPG+sfJsWyHqE6JaGTZ
r3Fu2h+wKGUvo/d5G/cDEBE2y7oqpht3vKfeyN+VtfB9ByMd3JDmiwwMP8lQMsLOpLoM+NH8qXXy
VHGU2keHb0Bn3nHEbW10+fjWkoJ6jeSP6S1Vo+L8Fq8ZJ1muOihzcexEOS+ecnL3hQTVw11ePcZ/
DZ/MC2h7bJf3bKeXLXNEyyQRZeuNuRL9ojh0UVst1rKrlmSe5STsUpXMJFEPOCEn0+R0xWW9GB7V
MVbGZnWUTtN743ttTvd4G6cx8LExqNthIYoydMs1m2HAw/VMNIt3938uIGLBvkQBhqE6gw6R5CYY
YrcHnS1wqYQt36Ef4fP/ZAF2G/ydJttCtTJRLAgCQmMzYlye0eBT88vOqvgU+VeJGRenwY4l8adN
l1qEGKOducafRafgsqyzSCNYl71/Z0zoF4MppVZyUkP4AuBd1cJaQRuK7mY8V+XjcH2DCH+6zdZY
gAzqC9oq7P/DeAXi3sJQpdBzoou4AiS052zgAgGSGL9TmA4OJLk9uhGtaHfQLPL57az2lRwYJCED
D1E31UJYWuG1K307JemDBPE4Ct6T8/TPsB4QYpGesyXSSh+3lbVXbsteycwCMVQdr7fCu8pXOnlq
NlYYpqlx7ZcX7MzQwraU3bS7NoA3zazoNMOSLL2hD0HR/8jZH1g/VflsD3pMnvypUtz4Qxax9/6l
MO3GinaNFVMZ6xl7WiDZuTP4w9Azowfzu0fIBZwgnmU58hdexu81pfKz4ipHWKzNPF87ui8oo1Xb
w37rHSRpnaXGkBygbrRXnEApnRS9Vpt3I50gBrqQrWUSI8wDn1g+V67AucyP1znDtZ0iZJppAg1k
wlz368Xodqzl8KUl00kDIG1Y9W/kCgMZgyEi7GA2NZgGw0IBi5M2ZcMT7Keqd26VUrVo3qa/eVRo
AzPcpGeJBakYMCkm64ZCLsqmkT0AImCO7/KiuMlWHQdOhk6LgQvS/ucOaZ9KoCV5eEsJ8WbhAc2D
qzAQSi6X7++45LtZybRkeAp8KdGNf4MKZwfJdpWA2AMTZgY8gXGri0mocH2Lxx+vca4I4xmd6onR
6VfG1Ox+hbgQ/5ak9dr0xBtJRxI0wT7OZiQgAAOzVk+up01wdHEneNnDAFn92CGCCgP8UCl10yXK
HQz83dAwz8K8JdkBl5RIqyeT6Trls3afgUiqB6bEBXd3fdVZsfNFKxZCqhMe2+lv6ew5W3/xZ+vz
NgTxQsoC/JJ/au5Hsln4K4TUd0nSVjt5nn6kQbNxzAXoxwMeZf+1M+CP2CTOX9GoNtt9crQ7n/7Z
7ENoeS6e8+DMcKSOidqLYJaUP5tAc7WP9CA22sFy/PVJbvTc/KW/bp0zZuTk+xRedEETVZV2AOGQ
BNCJ6+93vgrSjGX+e3TUKlKmqvwYw/UsLiOSRae+bRMqXOmkP0skbyULJbLO3hm2pbIvsnN7woUy
CdcAvZoalqXrXj8yAhtXI1Caj99x5NiRL74KqXuYw0tEaDE2FPKgANoXAIYeikHO9cw6cuzCRx8U
c8IkpgLfIQOtV2NK7lawpND/KR/IDuImpjsRYtAPMHB3BphJ6YMabfzJnlURQdPY8AeFy4J1FpCj
dLRmtj6xhJqhHHlWw4bZBE8JBJ72C2BcgdtG/6nnV8rXnxt+WvUsokO1xlzfRDZkmgG8lhXpxjye
/N1OdUItDcPmnOd89C96mUVNnIvvIp0ce0ZS31Ewa6LoYKuYKrTNvY773MEA7ME8axtuCH0tD9zl
5Uip4ZG0Oqg8IqEmh2GrzEu9aaAa2AqwvdWN/cpWQn0BKFm5JzIuY38NUG5rCXVC9wycKyE71ler
+D2oJKSF4ItOslpNvtoCi7u/M2aUBW2t92xDjfh1sbOwaqMXwM+guBOsusadRfi97jHsLQ8nj4jQ
Me1qe8b32sc2rCqOLDMnc0yDGYaj4YnpjNNTHTxw4eqgkT8ObQiC4ZbWBAeU+Bhz9IbclHDiXuM3
jw36ELFDvww8j++BvtSRzm7z6KDH/5baGBHncNlckvaWANmH1zEhD1CmZxm7va3wiRfz/c2C6zhF
o89lU34apK7QSfeBI5NjY2OM3NmtbEBRsIujKhPONashhS37+joLGcg1BZ/WgmRNmuL6HcHHzeDk
2rOeTcpVgF43rUCUNRzF+kszCMkGc70Mz70wEOMHKZo3KNhHnNIGBuxI3y0pZCAbeAeb09X2rqvf
GZUkyOy0kXUyu2+2DJnOksKHpkz+AlM2we2Sl9r+w0BeCoXxN3/J3dF8r/OV7npBZ6iN24nH+wlS
aLmwr4ezUu/Fwqf1kgoMOQTqTh5sHw5bM9Bram5pVpcdTr/x9cGaWvHQaN+WYmxov0bog9mhRKI9
ZmeYDmZqDwydjglGsWnbk6W0oCDZuCw0oKUeNdPCbn5KDxRyrGNXA57GI6yuf/X2fEWneR2EIZry
CGesnwMmuPB2NAEDuv80KdqK7PCmD4A2eFw//l4SyunNeNqCXSDAe4FuTIP6I5jHxjZPt5TL24RB
rcPbU4JoYSRPRJGlV1nv/apEaZI8d4IF87lgtllW+ZbnS5l+qakMjRI22Nc95JoYVhGt09ldUJzB
Stk6DGToMV2WNPu4HuQDCMtLyUfW/uvrMorAtreeQbyIMrRZrbOc8vntgVc8tre+/0pqYUAsQthg
pf/L6TMITXxgyaUigaTda6UTsQz7F6OQCS94ZM7syBZwG+38RBX1jw6kQqrA6zb2FehedvH3ZXa0
25Z8qh90aqESoBCTVXg5ohpbHIbSdO+Abwue8K92oKTW6ki+OA70lwlhXtFq8juD1XmhEtsq0o9J
0FU6tntc0tTzY4RUCUcfGW2phOqZHFIFrfhkUYjJfDCvC7Fs0y0qZEMmvn08LRFXY4c+NYGpijJu
R0pXpw9QgetWYTaEFpgYw8mrFqJFjvbJsHL2jcwtKbbI0lYDok1wEsUwM7eJjcZLcCFjzKsk7SHC
i/QYt1PSEMak+0mZUdzAoSCvT7l4o7qQnnlt98/KKoW060lC2HgfrrGjOrX/G23jJsrziHu13wLK
rFnBi1+CIgabo6j78v/JT6VKrk7kXhDycIVMhf+nIZIxIxRgltT1zML0DgGcB3nXto+gO5ZK1Uto
U/NA6yqKKqrL9sMsdvH3I0QrUgIUK12YSLyc+zG0+6bDFz/8065hsLlb1qTEnCahiRIW7dWSMHzt
uSNR0DW72lu+LBgnCBa0CL/9BsSbVTD4V7jctPXirTlzkj18uZ6qYVpq//C7HiKizd/2RGvGKMFM
6SH/LJBs3Fz+q0fa9BmZq2lj3J5MkHFYsxgKMaHJwcCHPsiI6k/h+qk75Allwg/hmBzB6h9iDqZo
6BYaTZht/et125byH7A4wMRHlDNYUslxXgNKt+iWNyiSrntJOIAZXMz64n57KAYuHDDP5Lo+//5O
cebH2AecWvGL2sG9pksMRE8soDVgaankRzT2sI1gjSHfWV34O9wRgYl8Uids3QHSMy+szEm6rlI1
fltcQHbZMRU1AaGedkeGCvowcq0ULci1Br6ikQydfctIhug7jPRYtc6Af9K2h8jKQSyOuVD9svt6
BArXo5dRz5cRJqgo67hM5kZU8RCNmLL2MQOEf0MrhR00v2cKjx/TVIlqxsPY2vFW35UKrphiPOba
xwae9256NEoTNfE8JLkfRUXQfqP4VIaoY0nsuwyOjlTRUTU5OsEWeCVswmFrRvWpbF2Q6G4EjuUS
RUpaykGpWHMx4u+NwbWBrquSKR1CHQHgXYFc79ifEjYfsKqYuP8sQg5vxRehBmekpxCtirkdI+/e
FU1ZJy36q6fottspoxrZSa+s3MH1w44s6QcKocxRvwyzTWPeN3yJQr80vd+nBINi+xI/b6II4WYz
NHsT3GASCj0HggAiOvm/Rsndn2H54tEXPS9wtSSNHucXZazFEYjuua2gKAQT124PrNcMXe02szoL
MRlMU1qpO1C+XwiOy0Uw4zCHec88ElDygGr27TckB1m/ui0mZ1uwXpqfGOCU9S+D20BnAH0MpPMz
sEV8ou5PBQOLc6TmIV2jXs8W2Aa7reTAmRT9Xe9dZTUL1Ho+FyljOcDMJ1N4D1W1JZJHFcdFbWGN
vywR1ymQvzFcuYnRxXkYeG5ZhV1NJYlUv14UfkiifL4EY1kaj3h7lrkqy7TPR4DuxXRdpOTdWaTI
y24rbnKRLw7dKlRgC042USP6/+FqpcPRr2if/EntKZ/zJSTE3GseNTL7H4/aldvBsfz8cxy4+Wuy
NOSk0bRhjDH+q/saRWnUDESe38UAeFpKZ/2YVWLeMMqTsiJO6kzZwe9ZW0XYTstmXEAHNKn4BpAr
16Yk24JNG+sX/+oRRyUtHmUQj+37QygXvLKbmw+0WIH+Eb7y4hyElx8GbtZuYHTjbsbaUqeDECWR
ZB/ENTVgcT72psM9RbyUGrOfnXMvEF61qBLImQF4M7pgSf/uyrD7CcnLWXGxqdWRPFKa+4Pq+JQo
gVADf41t9c7VgqtWfB8Q6wRW/wsywSyfeWoa8uK62Jx8I9pcoNjBK4UusdKBE9pk+Jm0t7V5wDUz
+XA6upYKnbPP2xR776sESacBp0afx/lV/IxiFEwA8vr+Zxze8C7d8goxsRKDwXbAz2QDiMkMHLxo
LFnp41v6+3y33yZ9lLid/L0TbWDLtdU0UE6pIwT16vsDPH5u519FFGFTZnFC+H4+M6IYFx/UcXGp
fgth5NMqxDdNRfbxTUG/yCmnG/BYI+c242vrv6djcQelFFlLAcAccFxJbZbuLvgm2AOj86nmhYrO
Ff4tu4Q3kx9AQhxQbgD5EJtkC/I4ETy4AqQSgO5Y7JwDA84LrVdN3/OAFSG9ygLElQbY2/oAoB3w
rzp9E9+6ww3bpxyVmdopMcKKIRnNLA8OT6A3LfUyiEhG7MPo/1f5HTPtfsA1N7owkIKMAvSDKfs5
vVcR89lQbv4gnHiFO66lf8FJOwpSlEZvJFArvsmB44WUtnGs7hd65TLcQ+EZIJqcGmGsruM4cGzs
sJRv0POzkJUYwntkaobcA2wAvhrAuJVIjUbX31E0RDFLbipCmzM9xDG2i/Iz/qwIRePvJoO5F684
C2Hv8KNoff7gjsqzbPcobe4TNNnwPFS3ByUH/0hPJnxzDm4nZ3HckaKm5FHEAnnKL9idFju023Rv
FZxPzN0SJfGPjNEkgnJwPdgFFZhR4GV/LUiOBhegsnSH2MEQfw/asXIeTxU1N9CDuhQ7TM4kJFI+
jnG//4USzU7aVrxvN3C/VFC5eLERw9XwVDyPxVoKyAH5hdZLGgPS6KUQo6yH95EP6ZRaetPH4bEf
BA409nvllV4eU8/kT5ENav8bvx8tuuM0OR1MM8hnd31Je2B9s9XiJnqz9dvIAVLGrbSnV7330Zme
ve5ZaI5w6VyG3kQsOBE1VN/Artsb+Tsi7yb2oeTPD3QhTFvqBU8hi8gxjs3GjM9r9Nf3ipw+rVOx
mqeGTFDA4rVnxEBh4l4kUWY2PcrPRs9X/jEXCd0gjM86lIVEA+eV8r+F9KTBsVUuLdjVyFU024ag
K2ET34pmHXXu0SFWMAFrGZlFhSWNc4PBiptIXl42B/PNQBHiESXkIF1qL7atpNujzp9csed1hzkr
DGMa5uKq8Bv94zIA5/f2r0E4P4f/32nGN9GTqxge73c+tLs0FPyX32lbok8pjAR685aU/gNBo7HV
ko0MsUwuUXNeDWgqeIP8bPt1rY4bHkcmaDr7il5ydYSFgqvew/KPa8lZ+bcG3EhyxqpT3wqMD6qC
Z46perazdIetdNdwtUGTzj4NVAlbJbFVDWX1gdY3q40N7iTuwsy6I43J2BheAcc2MqlPKwohgiAC
+TypcoHTM4mvUeluOx18R6r432C1psIJuGuONPU60l2xWKFXQduOJcIxED8BWnFzgbkDuCGaJCe7
5sJAFwsHyZTFqH4i1JIqsIq5fr+RQ4Zb3HZVFFq4k2X625hbrH+AZctMlOPZbqL3kSAL0nFgSmvQ
745U2UiYYCppjaNqci8BuK/gG8xX4gkyQ0TJiCn4NMB1v9+8sy4pMk0emvidPvNOL4VscWfmFwiL
nEVNCTrRyYO9BhBZA8htFrZ98BiP1B1j4yx+evpNAT/1pUp22FGlziSAIBHVBj6X0Yj6GwsYPRN8
aLfYzlrXzCdNpU3TU7iFBV3oqx/QQ3tPRgkPx2v9tu2LhwiaFNLVpUNkCdAZLuzcLMSFCvkQl51W
kWOTi/8pQmq5AfDwreQY2j6G39FfVVItSnVarEVdJvmOl1r5gaLPOBs3Sb/dnZ23V5+pTmQRd5wz
8dos414j+rk832WSBDFpGU3vfo1kKqwfFH8HATYTW/3RgubmMqLtCR+V3EA/ruch/bIDeFKZg2L8
SfMEqREMS/mHiHuafKGMd0HSw0AB3oif0e+vT+BczGywCE3n7tKT9cPj6dzKvHBp4TvZr0FbaXIh
QHAYUtl/eMhOJGbvVJR8M0tQ+Dv7lXi7g8A6ZZ6gBSGebpkRinzGCPhm4dkF+FFdugutD3W+7A7U
9GhgOcwahNJt0yb61TuN+qV+7NuPi1C2oNZsASrp+R4hro/vRvIkJiIn+iXpYBV2em9Ne3q9mYcL
vbI72CqUrZJ8aCIr5cSNNEYt9yazXND+WOZwoQl2/3ANmdbns/I/UCbzFMLcbV6ZDIhoFc3XyaS3
2sJ+g8PzwDa8rTTJmWR/P5X3H1/EQ2M3il230eSHJcRMmkWlBo3XmsQfIIQAAWf5GjdJNgcQxuu7
82IMVWF2AHF7vfHqAbhiQELs7dCPqePmOBxR5jNVsfTfl6n/gWIsPPkxz2BoSR0Pc55wvhLPKNyQ
8oRTqW8y/hhU6TeOyhe+WpxjMAay+OVikApdVz5mcamb3ueg734eX6hpuLWlv9bOWUDhzlOn88H/
MlqVcRIx+jw46v2KMS+Kr7hZnyW9HMrRucWtE8HbZm7HrMkH91Y1onHd8LubAcIy51m//StqJpti
ztz48+cZC/FGPXBfqoV0ttwCSTD8AABG2Lc+/kbANzHsgBE5xkk8YvcdZbFg/oWJuKsB1y0gCtYY
0PNIaoKsjzEVUEtrs+mhCyuycS8InWQrt0rxfq2ZNzdFyQ8H+8KUXUPFg5/p1BeKQSakSZphMbsz
/DLHuhMwob4WBDefU0TP0Pe+ohrKGyI9nKv4lU9i3+/LqTxaHctyHHv1HZN+05YxJc0+tZIBbHub
PsTVtAjCQhy+/3xBn/vrIbW11G2PEwtWzz3RW9Zwt1e0bZzZ/unLLvn9tfp7vozXoQSCR4PUklrj
DJxGvwXUIldtulr6OoJp8qzMHhXXNqik/HNGqGxeZaAx6PoRz1XZVzSo0YqdqGvC6cGcFtjPDpzM
w0u77EHVVEdAbA8ArvhqCWunrkEC81aEo8Ud4yR7Fw9XdnXHKEqiO2ybRiqYjYy2hrnnqjaQjciw
M6ljsKblnxEjnUP+6l6/TFoFVij8Dz+h1bL77aL3AooJMf1FKJOC6FiMu94ut7UGFncTNeQZXNF7
LcT8nUmhgofauzYQ+LWDiRexypECpn0dGugkOSSr1DnY7+Bqa60nPqv/EDq7UfT85tX3WViiJXYL
6/MjSqpKXM1bw9aJycKvQPsoQuImT5eodHU4P7l5jlcyWVYNqUIkPqHmpOlPj+mHQwLLbMxTjYso
KlTV04mvS5nAP2k2SXq7xGtTR7mWzkmFsW1FQwce2g7tD2BvHtWkiwXpEkRvIvegznAm8HabrwX5
EPa01h0gg+4rxU+53LIWuReJtTf884V1Iu4JNaCSqum4d7MWI5osBLimI6tN9l/axHHFjuwuud4j
JbzAMGiOAGYZlvbh0muN8VZtfg2VMz+fjJ0ZCMQt2XNlllm/lIiP2iZXdCK4RlgK+Cu3/QTsxWs0
8ShAGHm2R5rYEoCKmqYctYtNXWAhUnMMz+3yguribikEjHFArNasVgMZ0gUQGeyc7CIcdhiEuXdg
4pA9MTXw30oruSwTgTRZLYBORteR0meQZadOFvcynUMXFvSVZc8cPuFU3J1jB9V5/h3vQw7D/F/L
MkW5A+osqmBqM4bIzg7yyQ+hmi7JWleoOd3X5k4LonIwGdw8lGhqd4HkE0XvGpUjObwnE5679MFz
fpUYAqQ4IjMgAvb4Foqpc0V6xKbxW2qg2JvyI4OU90FkKBYAA1jGjfW+q64tds4YgMiYmQgfCBhU
XaaCoaWQVyChH4PZqahOwa6x1tyt8F6JL8P5JqB3f1uB11SaFFudK10vYSurLRQK00seM+n+qQNB
XsMJi8kCupTEJbL6IxtNM8P98u4mU76WAl1X0jHjc8DGbL4TN7FC5NAz2lB6KoAyxaJwucdD9wGN
YEjmep3wqBPlQY/r+9BjGVkxn+n2c+ovO+atJMlQYCrr4vrbEMjUJzfsbPcsmYZZ/4AqBNAsrkZm
lvw00QS26KHbcYwufBW86HFCzkUamYBTpHXGaUCooOjy6EzuR+cQE6HOYldzNyQrXf5yAv8C1yVa
KzvMot9yhKg1YXzlqP2y1dGtuoDiYYTxBHoGzzQt9ASpAV7N/XKDmtkcHKOADqUJHtzEt8kJWat+
SYG09YyVfjeKqafAd7i8hY87btxTrJT1eu5fmMFUgNTqEZ8PYhaNELf0K/XvVWYVhRR5+mC/6gm4
2+X9OXzd0zdYmyt7HgGil0gnTcLmLVqj2Vs0FQGdroqTMCWERFFJOJzyYyTHz0uweKILxE2uMVex
Wlx26mcjFuqqCGJO6r+g6/TCZpNTaJlx9Coj3XenKXstM4YNr1R1Jv7Gjj9o7t9OfGaTHqOZO9Mb
X+OXqaIhFHKEESrSpcPReEjSwPjatfITdg2Pua6O/8vQCCyPhUbRtwxZlORtv69n21WYQwOBqMh2
1uWukPpbfDxQFTnf+rqADVG6BOO7wyDmUbwHB0NCtviO5AUW2YqcRxg2RbutFbXGBGj55jUaTZIv
IPocGIwiXOnzlc+sVwZOheGq+F/S8YlqMl30J5/DkoJhTcpjGqJI+hr8mLU9WUVHfT9LgqrKuwv7
OUslLcuoDzkLdkTbvV3eH2bbMeyZO3fKu+AN6yWVoN9e6T8Z1XqHYzAsvYQjRH4Zp+bCTYuMssru
AJMA8CzaTXhP5fz28dJI8pvbuLjiHungEvw1ZMyeHO+NUg7dl8LFQmuuYz7lvLLbrj3fPFRcEWh0
1Qr+bzjHu64HiKGpYWL6oDbR9dC1SHjxt0bkCYTBJQURXbYAv0oVPOHa2gAEmufFaEromLVA/g8o
9aioarpYSMv1cPgOYlgQvXnNG0yptvH98k8R/M+a2+NQuw9w59xpXwyVgK1wA5ObnVxhXxHEXXmj
1Vt0IA9OS8KJEl+dDz+eAihn3nVnN9dpizr4e3fUM1ynAGo7xI2KT+Rv3RkfI7i34xygA2dwqKsS
R8x1IQ31crV4c5YR6pRFA6bJzOHUN2+UWN6I6lhKpTjuV+4Dr04k2uSICCvKYvBNXyqltSo7H+TV
zBgPDYqYuuowHGVnOrxVjuoPH+R6D4jz4NAJV00HvoGB1GkpSEafx39aZq7lz0R+4SK2vOfOqvSB
YDyrbAST4pVNP+PJ/UylA8n6QVjHx39Kt/ViM5lnKr6TGRUqlrHBVaSF0aqkv6b6aBhHfdeKwX9C
lTDFAqfdclOSrsQgFoW+ZwkRLmxukAIiawWU39DMg130vY6Ub/kPrnm4isCXhhzpa8tK+stah1So
DIQQEJh4A8WEriH28ok+ORVkB3DvgAYZa2TPhTgQWu9OhhP9BpH1Cmz3atZoQLPhRFTQ0sUZra4a
DztrANgM76kNclXRBv6dEuN0ShgSZFshYOHQ5n1n1jmy6ESskjT7O6rm/uWlgpoTyG7WU0tyXClS
ngVjNpbIH+vv6lgJXIU7oGfiuZ5L2XxQ58ivx2FlkbBH/jxNAeZrLgGyg9E6nQDCZO5ZlgcW3920
XRdel6b/f3YsUznRQcw+ynYG0XAaPg9mJQtxYQE0cy4EeK/Y8QRS60wLCNxyTtEjz0LFvrvJiodv
W/Knl1T9S0f6bGIISD/NrPHH3DL1N2AqvKU2FhRXrO3Uu0FisGvMrKRt9Kv79Sg/JvvphVL2wckA
1O1kZN/zymxVGruaaRgBbXFwaNsEGpaW7DRfgYZ26GXJtYdm/R1+9FTj8+7MROBCWTMRKecsL3ux
bhytFW2q5vpv+GVLamDUQiNpQEPMoEwx91wZDCUZxucDIJ9DCgCHqcwOXR7e5uB+v6NtQ7t4zJr1
SBzH7+zJm0MO3tuw24q2nG2l5G0WJTWQOpT9oPDFNTdy0k5522rsti7ewgAbeCgmGC3/criyo5Jz
JF5Y4oeRtohd/8wIw0o4V4V267S5juK/4b+0SszKf5YQa3Ioz3NqtD2JHDjOWLJEe+9DA+LERtEI
NvAvWgXgWKLIPF2BXdnw+mzwSpBAsK/311r8h4iq3MgqKORJ6m8bUFV3CJrU5RgsiRtKA+ytugK+
b6MaRBxTCkpa/gd6agTtIr5sxNcIroTr36O+dsSAIbUyNlD3L/vXS2i5vABSML3JgyNUMByNPLrG
YBzTVYOjQ/zMsnso2+Fdqn815+stTDhDcwYTHyIjsdv1kzpW6U8qCiYYwmObHdtMWp+QWTx/2Pgb
fB6z8pigFXVk/XMoRcrX6CEDz1RwHE55ypNiGgtzJEH8vv0bO8OHdD9cZvsJX32EB1ffyxW0JU0B
IzhmHRVWG3a79inkAdMEVyd442GqmVq+SCXKlLq40VCs6VAoPWB7YFKsp0yVfKc7IQJgess/L4Mx
Kw6tcJ6I1OuLpvxrGlMnsX0Z63syrlHoF9lgxdACfUoQK9HR9j+tbb2msiazOZ5V/rW5gtJfKHlo
hwjKK1wqYI4wxLGW7EAu3SuIWuIZShFzr1fQByZe1GtAA+WHiMYpfftcrT7kfc1IVQFIf3PPqQw4
NpZC78qrmTiMRR3BI/vrXPXEVlmXj/4r2YLj808lR8See3uwP75TOPRW6RHm6kzVQ9z8iTbheCHc
l/EomW8G52/l4k9dk5P8LYtiBtcEXG28hJZzaTbD2DESceyxcatlUM8E/7eVgeyaxNRLkJZ3faEp
atkc1Bdtq4xGZMD7ATki8fNHSPV2qtFEChpaWRosJQ7of9m8VQfn+/slOcAZ4DRgR7RbQs1psP2W
GCDMp186h1aHOhVY+Rz9SaU0v11uQnujVemxWQZ17BIc1kyYTO2AZAhsUiLhUsVs2D/W/9IPeDkZ
nJvaTc1UZfkM88KNMkzkX3Ah86Wl1WK+BI31yvkIy3NVGUEh/PWYioV5m/Tq3LaxNJZ1AAJKfp47
oQxwlAKgId5XjBQcZldf5s7H6W6VIR0jXNwtZ2h60/48OqWBMt6OL5W0fEhUhNhsL9l9dK/KCP9L
Q8Wq+vIzYBj2so9RpUfyHxEQhHGVzWRFxa4jnCQwmoEJd5KdH3yaDdwdcF8o0HGda4T5weVxmXnr
6j0cBj2dtJ+8OSW0obif4rmFd+GJcBtR8oxLrohJQ6A6qJ10r1meDGCsutcYs7PtnY9o842Gmy8B
V2Zuz0q1fGNEZvx75UoHOI7AByRWOGfce2mLUziLOnQjr7RmYTkwZx03LnCk9UhkVgjs7+63KFVn
VZsbTBOMAE0zVJmTT/uDh/w7GglZLMZbdH9ynsH9zP8Y3O+5t89MJ4LdBNKw4As3UNU2OQPVPrMT
QKTlRv+CifDsmYYPMPRWOsL3qooWec9w0/cyEN4/H3/jHrruL3a/l1pTh4r938bzd8bW1/NebdR4
BuRr0G/G6wt5mSo5jkvwOiXduYxFLX5S7NSqwIGsnEALdY2p6e7uzkN8Vjsz7EuG1mFc/a1lYgIR
KhL9VUPUC1BkZN9X4QoJ9E216p3UHPtsEQIXbLo/Agw6Ehq2rvuVCpYmlEMpWJq7Ld6ETrQRGotx
NSJuWrARBh2TDx20lZePVJjPvstp6a9kJDl8vnwWZkcgALo+NUmKbdN+yMecuDqITdRYwqO/hdFa
BYXDgAxGqA84wUE6h7HHRbB19fpsL0ddrU80KNZUrrnQRt7+z1N1OV23mrKNrjT1WLUQZsNwXTi1
4tAuz9l3dudXiG0ZFy5VWqyJaPXYMdhE9vKgjrG760tnIrivf47+ZSsuwuWErBldLnZTR7706d0C
tHz6y5w1Q5Pg3HbS/FxPJNH6g3yOntPaZcuus0b42WkiH09ccBvyRD153YwdoNI3Z8Yad+FNkUcZ
xwZnwVHdKAgSxt5PtGplupt8/cKh+u/tyiQ99GbUm/5VSb8Gn3G2dExqHfWnG/FFzd+KPW2vRTiN
W8APxxeq3kl14QBv7WYPZXA/S0D1fnRNKXowG4zT+eEVzs+nqvUJxALsxg3X3D/ttnJMs/vMLbHG
/Iu/35fnbNCw22M8r0xF9r/qDZKHqtdyKmpe0LZOtlrY4YbwIg2GoTSlD2y0gdenOL/W5iwPXHWd
wj+W5GV6Szu+5z+ctxPNcxtzv3iOC/Id7Pu7v18T/VhLAEEiH/PyxBOmbfPS2XbgOCmkBmVfoLQW
A4XZrL7EDo7jjWsuL2wiiISEBYoXL2t/iJK0h3aCcg63TT6piMGBbFHlLIfyH0KkfqP6Yh2cAILH
iSzSbZ2EcoauRZ6ti/jh0+OJZVaUjS2SJMsAi+OPJHC4MIGUX+cXdr7mh7SCOy2shxS6mYwiO2a0
cqjhjLxsDakk5AIuzfTVMtddiIghapH7zJ8hjNNh+qYhFWEGrNy0fJBJ2Y4mKLYo34YSpzSR7H3F
+LaxoYkxvDYR+oqCf/UOXOY/ECwSY/j5sZBGmNpTKXMAb+xi2n9nmXxC0LLmueaybzbBOrhsdjh3
zVibQ2LMMnGtSKNwU4KfUyYXbT0gr+RAn5dRBSHblTrGJUl+t9o/WgL5JoejKWhSc02q0I8roM4v
KmLEotZPSWmbfl5Pui5b/plBqsvH3R8RNu79UdGPcXqDKIdNTongFt/w9je61/NnyDcvabSMQKYE
L1rkd4APepA8qLAp5gAHPosrjmLMlAs6JfCkkP4hPiU6ZblU856M/0g+2IsiuJMJkH9RqVlxNuZB
d9BhuiaiXkIeTJBZElNtsPN0Fk0fCLufUYIQ4uV9SxJ4rVd3dgFc6s6VMzm4v+rUDTJenKBzTEOg
ti66JC+TzvYq6Nspf5Gd3VMzsSlFmG0H7LnlMrIT2EpUXPUHiDLcpMbvtQ8ScPTNaQ9qHCROay4i
9W5xhFiyClWiwlhAas3vFQRm0luMtUpjmU/jFuDFdIJng9sENlPjz/NXHnaGoRrgaehGnoiLGcG4
YsxUMQlfnj4UNodChJd7YU+dHP6HM459TD8a3AtRQRfWdNlnVc7E0BqxEJ9ZHYV43r6Egezy4XL1
hr0lLnslApGFLVNed5KPMjPEE5Ez8F1jXy4JvfgFpNS30JaN2Ux22VUQc7BTY3m8HmsUfzB/gpto
ASZoqdaEObWelx4LFmMOFISMLSVyCa5uxBDGs5pA2ZI8WERTM6qK179JJlQ5IxUVmpf7GW3noIAu
3Uiz36TYt8og5c7e7TL/bz9NP3Lb0IFviT5AbQxrHU9GQrZLjrQpxasZi9kcB5SZswzzgqJLeBN+
3CQ6rIOTU0CpKnoF0CRO56D64tL9pts+d9uiciGuHuJzEyQzaH/U5ybFTJD1PuTcpIK7oZsRrv7W
WORb81imI8vKxHitZ9sKEQQjPZ1pJrZal533tda5BRlhprpz4k706uF5pKXAdN9hj5DPId9SSlRF
CkcVTSX4RPixmJLW3m1AEbUvIjxL5L6cVIclr00n+9aTZQm02mwYn9UBY1xRQgFsN5foAprUYPHT
rKJ25qCBHKarYcWbdvVD2Vsj7QK5hGGVYgk2x5JNnaQ5iDg2M5EOa7iTAGDxLONNlUNdkpahlGss
546/e2R9HrLjRXDXAwGOo6arKfG+/p2CuYhavxWKw8epw84Yunh1RPnr8sRud+Z1HdgTMWWi1i98
Ktwpj1KoyrHaKubFEaka+kbdNuq4pkSrN0k2jN+KymfLr7sHBhI3qOzSJrcgggaxekNRHIuZRrQr
OGK+dBT6yLHOrw4ptwZbn1407wcYD7ifKVyRxSidR1MJI5dIyjefqj8NWi710FVxckZuDdLPRpKr
lmlZ2SM86RNGD5ku5yOPQBSLRT9Q7BugnX7tLN2yHlAhUwNO3g43e6zLVC2mFSrqtcVg9feL9Ps1
YsffzAp2BnkrJUjdpua19YIuddkft8DKXfk8xQxANOhlzjn8gp9aRGKXK+ufRY1Ksm67RUnOgWaH
5ggcd3hF6FeCY/maMTSTSd75R/xIXihS4l75WTT9m0Jjk46WKb7KoKi+0gvvhKf+pBEt7qDzZj3s
Rr1llSGwC6sxNgvzEZDe+VBuod7Vfty2QqVuT4exqFoI/bb0YyULxdEb9yYmucteYAOGDuUsUSjP
N9mAYkM9Q7Pv8jC8EF/6XX/oR1NQXav8+bhGmnOpdasTRDJfoWyUgX+AosOIpV+LiomURvWqq/uT
g4w9u8crgYcHIxZEpXYg1Kb/91+K3Z5zOqJgEdXp1ptFpbWTSL/M6HLLyde+XAWvBDyIco2gZTvE
zCtqSxyBwxSFKQtbs5TPxTQE2IP0aEERTM9Ga14URkVLzQM4GcHjGzYsbVGlXyn0ZW0WIyvaqGVx
FJwBgq5KIjXm9SF7/sWA8UAxtzMdiUIaklePKPuplciIk4J8VWxeCnETv6yFL3S3DcC30QOlLB2o
7x4nV/xMZaGKr6nRS9sM6Ls28gyRgw8ZG9LaEtOjvApJTSRTySkbEM9dj28OuTx4XcJRrRFIve/B
bhpvJqfqIF/x140Xnr13Klcp9ItuoFeflnIpzV0xFI8LxDpgxvppvRkdKkuKEVpZq6dLVEFIEahi
U4T/YzhhkaWeBtgcaUR8N4xZLHPt8D3kEA3Jsg4qfyqFqntzqAujOB9zo5rWJ0vMBl93g5Ih4y/w
jj8o4JNDS4j/tYbBPwUZfCgxaoLKSIwqeHy3HkP3IzIOSLp6wonYejgdRzD4st4v8Usl+NgkrtWF
0Msz8J+SS7mvv8KTCxsNYJDbgfjly8LHY1A5cV1/PpAnqa8zSyXS9ZQV86uw3A8mzu2NYMt85imQ
ev+xOHc6tI8tSxfOtkMbnXkiKB9+sPAy4iyDeYp40L4yqSyMk8SZ+lNTEE336lKOvsXU8oNdgY/L
Rk2OHC8iW0ZsiRdOgj2JbX8Bg6yU9h2J/i45nxzuVTjYOxUddYuzEabagwv4RMw478dwdDkdjRjd
7Z0JBRNmZyF2Wbyf2SI89efJd0hYJ5Asl0Dn0OQoRBoysGKW3b+DKz5Vmo0LsTCYtRk5UTjYR8+o
TqiwnKbWiuYrKQztFKHFRCSvk8gNxwfcQsGPvE5ZCRCAgi9Wzx370xhO8O0t/s44I7hddLNCntKh
Otd+ONf5lK5cpelV2FNm09ZEJtTf8T7jKqlv/rROdxzTxJCtSui4PV+nMkmCWjFjDXj4itFN4ft2
g9ayDyt9i7/LT76SRYbxYai4hU2i9/vD2VzYqzCdX4+FpwuP2DwR9IdPtk6DPDDtwM2kNpv+m3kq
ERXhL4vHvOvzkaxl41OxGEUZFQz20p4NVAPbyhhZCGiUvKtVkwff1flzKr2G/hJs/KbtvO0eE7Sq
WpOldzgGo+HA4aSkij5XMkaOnnh3qXs1RZN0e561RpYsL5gWv/ObC23lnGyFkW0n8jse0UbnCpGl
BXibMgri1BKNxhQeG3arRxqsK0EuZAwL3vPY2XplKvf0VCjztnFpAanBlVfbT4CK+n2/0vUhV7v3
2Lz+T7okfDZwyp0B+oL3OcWLqR0lgBH+0kxJxMhpxObdBKdCwE3w1f9lgx9LfEsoVvPnsadHMVEH
OaAebt1jt94+TJFgElv8X9LIRsATLww4tVQTpQZ7M0JHzmvdH0TofivPH0MgrehErUng4+L+xZCx
/yYng32sGF2+xxMEcYJsxkkvngZg8Ixf6WDRixdIecGrHXlw+JR1n7s5Uj/Kqxu4cLqA6Tw7/qZu
uRMiEfVJ+x+2kWIa1jUIIzaWoIsKWdkF2TPLKe/U1wKZHaNGCPSyHO54Y/q9vetsep45Z+zBNqha
VOkTW0sr89ETXWCAFjDdFcs0Vazr5yrrJKcD55/H5B+CK+VT6KVi0ACy91FqA1SlAjheE38VjzWt
UQpAletB76f+G+xM+DhldHbPmQ7L5c/3MUHNVdl5hEfoUpA0D/XpnB5g5nVdVUq1+GOJnfdUNQt/
YyG8GiyOTx6lKjTpfRBTU056VXCXHGtSbGVdOMBNbXjRMHE9j3mPsbRt1PTQbvHYAsoFlK9egPo0
/FjNsSacCbdDk7opWiNs5J5bI9MtTbttdiiJV56fjEU6MrUcvydhekCGpiNPvFDNJlJd18yxsadx
w4Q8SXfOh34ey1hq/O9MSl/M23sO/b4YYQySf1KVOpG8u3DUsE1sBrzyUg50aG2lfKJX81WiRHjG
wZYC29XOGVZEW9Iav1cX4tgbYfNX8M3zX7E4/DJl942obh45UyQDAlqi26xWZ4hlzhPlLlqQ1FI8
KjJRhJ7Tzh3vUfxH+iRNfsC8u85vOOuh/EK5mUesRG9ad/PvGd0yFb3e/+08sq69+/zpXk3UR7DM
CrAdDt9tN8O6CRhfl8RqUqYn379yFBsn2fckDHcP01h8eOF8EfdyRQoCGfZnWlhbVsqlLb3gBGAI
nN28V+kghwfpR7p3+Gx+bGbzh9qaALvwtpp/O/JcyxEzqAHyqowkCCH1Yl5olPYhSwkq7qFTmrul
mEJREqMIhCshXBzPdSeTAbGA6ZCsdL9L/o5VMwAFLDmGGcCQkEbDbyy0VIu7clkbfjtHyeRMKMDx
0+7ajFKcKzEp/ve5xmsdGZvYpgc8VSUn7IcleyE7oYXwxnNKfrRXYHEBRUsicxl2zWbypdrnJegI
0QmQU/u/ut+lCpRy/4Alm7QQ3rqUEIBacLXM3Fk3yf3ssfKL9ADj974PN5lqbJ1kQJO0QrzSIaUh
DZI93QVRiBF7bk7HDQOAkV+eBy8Nk78Lr0ob95Ee0E/dnfpqOVBrxS3h9xjW4K+3UraRsBVPeSLh
NR8zTzcXn51zkJ/dFrQ6+6kTsb9eFnwJ+l0sCryLWvohb4T5oemANXwvJx8LVDZZFK44DT4ldfzo
AjJk//DJvP5snF4r2cx6Bs0P9k5fRWaHdp6NliUfJL8yxVhaqVPsXS1ghykz8QKjaJ/qCnF8d1a/
SxSI73DzVwNpj99DZXF/aN62BZUvBNf1wCTSl/JdzdWodMyPaiReyiGmfe2sIJv/IKJ3f5lOnVQl
zenUpkrzwRjtWraRKZ80eN4z51zlBRL5tS11KEpyGrj0F1OF9sSv1wtJ2UK3oSyR/Qt3JQ7DFZ5e
b18jqogCozxW+7qbJnAvAL5dnO3C/b2LdZ60gZRvcMPFtnR2wgg/gJz9zbBwxDgWY4ACX8yJp59M
QnklhWDIT2oorFDYpV3E+QCQ41D66JIV+6oCQaHWMUqc6uqjqxK1OoX5n0S5L1XNEe4+MnNoQAeU
375q61l5JkdfX9oA/zheOXBwv0ztHTNEKCfiEwdrA7HEgnLmYRL08VPzBmwNuvMXSHPDys8MQvLF
GPBKS8WNe3qPXHzSDifSX89AJXRIHGlArpjgCHelh8f+i8eG2+Lysj+JXakTROaoPQcy7MaKkBRb
1yYaEcrNsOjU7pmJMvuosLmM2NGfnz1VdVaKGVVlXVefrB4mI3TMwcYKWJH/TlgjYK+ATn5lJXf7
MuNOBE7Ebhn8U/NHbgvIMItfwGVOLtH0sswssDRzq8YA9bfRVEzuNLMnEivA6RfgOcSUScQMMd0j
oNA5XhHLl1ZqPJDjpFOtoplHlpl4PXqk0lqkP+W8cRfLKm+8a1PAbBSVd1/8+gfvh26zpFpA10Je
owkW/kh50Qw2h563mjB9zHNGHWJe2ZvvcwjHOjiX79b16GIFG9nuGOpW9BhUVHZYbufq7pHocffi
3IwljLkkc9wHD+dIfjWmkBfxQrRS9k1n0sWVDPQQK6YZ2d+VDVZ9d5rYwtqBz6PdGTl1w+ouI5OU
PN0Vu9xazf3amu/O3BK+YlYMYozgkiSqGOC0RRyy497id8MenMXPZQaWv0eNWkaTPdKveP9+JsVe
/c1lVZEIYPiQ/f4vxpDDTTjVKfEBx1cdjWreWuwMQOvio7L3/mni/tAwQ20J0cH5/h0ODIQpPa9y
wqlpPK83OdlcKZRxdTrJdMmGo/qvHntcorGRk1vyxIGEL9O15yUtOtwGi3pNUNfxGsy+QEBJa12w
1lZxE+0Iyn33I92IUUQsbaroTiU+L6TiE1ToBty1wxM62Ep89YqKl7RLDLrjo8wc4oPfkyULF3Ot
TQ8VoTdZltRxN9tUlMtqAtuaQeF4aYXpHhu/RTC4p79lCjRL/l/+deNlooLq1uVFvM1QSkkyWj9S
hF4dzrFpKwFZVMK2bZBj18XpqXFhOSWGpedAwGONZfE6Z6B9fwXGwVuATwnodrhXvgC1h7ym2et1
ZL89muA/2UAibXCvF8bMpJglFe/sQYmn0mjFZ8v751E5ykN4uiuTiRVZhbM60WAoAmfv60q1z2Pq
dYvasI07fIULmkRX5g6gJTWE1c9QiPDbiHakqy4lR1M085+8LaZLuDXfZVYyjnu5CjRtpPLQAMkg
cjocgia7yS0JCE159tk2AfCwma9SMBoK5DGJYv7i4w7IteaQUgiGKwJ5m72jIx/Tmv2zb/E53r/B
4kgy1lzBtuG1j9Mo5qhIoinjAKb4OjZCRrWS3KINlxvjYY2idFNDy0RE6dYhCat596SXaXKCw4Xy
nzf80yWEE/+ixc/tBSZZrHsmEJckWhf68ck4cepDAHYhaMZVqiHVgtSSMM47dpubVl46RngVnG+B
Rp49FHqRJX/hBXIbMDV6NsRmoReP1a3Z4hzIBMgcooZ/HS1SZ+PiZX/GAUI+wl+2qnjW91MHLE1Z
e9EeF2fmV1XQ3yV9vj9AoiFoxihRTylrJLRmMf+0cJz4BnpfX3OCfHetKg7hbTZTQcCaxYM1O3/6
FYyxgY/qaAde5o8lAiOMrWrM+sp1KAVmgCCWRxxoKuh/0sDsidGesGHUDu51OCwKEStGAdwbNomN
AP62jQWTUzITuThvOiFzYemX2YfRy+c3z0517Wkcu/Eup1qi2EWe5C9nt8mn+DzjTAaGflUAMJGp
EQXcrouGa6toCbSabp2uLzYH70g89aahd62Gz9zIxz/fG/dHG9YE0Dpvyhztz6l0sV4edOPGC0Ht
DAAEDR7VYjUF1+Ibc/Yn8H3N8KSu1tXqFn+MtSGZG/VR93XAlZ+PpSVltOcmBTbUw+2lg0sEmGR5
JlEF7dFpAXghHITptabDccnpk/4CgGmRwE9sjq1aMaoAI/sCiKJyVZeVtXfiBOsiK5JWCJ3lQDKg
Llo64EzeMrVB9Ha7PYd9isU06YGxOTiaamGEPlKJKsrj57Ab/82ZWfbYAXIGeOkGOTp6iJJo1nsa
MwkMZcre2S7PbFkEx/B8ZVH2foZ1gYqQNj6EpVWydr4GofIIQNCtQD25dWpJlzajPfpSFR0LVLJI
G+4cNTWYEQcHu29E+tJ1x+MhPO401McrJhuEUN85ot8mLA9MVVANECFYPWLuorSmKk+EYJ3qcl2T
PYwnWq5UePsTU4jobar7+bE433E7IVARplSx39F9lcGFtylr/DSauIf21x/vSjd29HG2FeVjHYtn
Rl9RH8d9uKX51BT0mXxTShzxX7+fuQL83a8jRIBaYwNYWzrsGGE1IGuAhO6mhEHCgoiuZrSdFe9Z
KV9EnfYBgkQRCMg4jSQOBhY7cD2RFXr7NLcJa5T7DLfhayFlTZhi7UP2Svo+b0H13Cw0KWHVQHcZ
8BRKkVE4Jgis46Rve1wFl/TArmz7HZLLfKuxiHcqEk1zOaZMHUzWpcfbrixhLWzW4VCGFX56Elr9
ldPQNw4YHDydXkTvsErDZToop9Ug9LdqjcIG5UvEggs6qz5fQWTAKBTafW8/A1TS7n1nPEhzRXR5
DFcU8Qx3L+VmrqwzgrK3TFfcIr2AMYesPOjq9mTfrvE+yXbFRX1NKmsdTATKQu6I6klmlrltjen5
1Lfktjl987/mzIF2A/ejudCTCzMx7odnm9cWgFlNjcrU8F9LBAj8jV1cOXKbx28CB8TpQeVNiHhv
/g+MTRYKBOrTjzlJ2tMyrCIiwLJ0FYo8nTzcjDbt2pWhaWyUTBBmnsHGaF4TgAv7CycbD9XcAMoG
FIZ7Mb6GGeQykVS4rokeHMiPm8nhsacw67jR6AO1zPARIK26mEsK5dRJNqhjVwxraPI72JCsIXOm
ZWRhfDwWb6zB8bReZhfWkIup/u2X5jvnan5u/cLL7GA/IXmnzjY8pIHzIqQmt18DukAFgX6gNpbd
fE4GOvjusrD2g95ALHRLs3Bfi3zKTqtOa9or/hOJhzGzY5BitAJ9ScKBtpAeKlTUmWg7WxCwB8eT
DFG+7w/IjXuU+d5uW1YhhxNbwF1z/MgLJL3u817yDCtenw9B9NZ42gI5OJO1gTSrmYD+jSu0Wp17
Lt6sN8UZF5ylPsv+alRJRrhy+Np8uooKa5L6mGcYkKUUFnZpYTSPA2G9eULiXxi1OvWY/LRmz2FP
oznPH+rpzbPC3i1PCgBAvucu6h5zu/vTZoQBUOV0hrbpmFjyfQDFWw0Hf7XTQgZVCFgvBkdJ6r18
/pOeb31z5NK8pwerjZfwa2rco28J+OnQjZTLcVbx+SlkzYf6OvUWNzR74UlAxyWbBp7mVc8vfWMY
vpstCXCi50PKUZFU5Gymclq+5MV6ViXnQHjDWoYXdFX3FB9RKa2RZBca1wyoWisqaqyH+efIMXwa
0eiJOQWg081zfhl2ZIHZaUUAy3XMIPocFdc+CGX82CXpwcReBFURzcYnqNAg016btM+SMHE5LoDF
AG35jdCNoXp0uefSQY8QZQwsN4gIwQyOzWuW9ZyPc7yw32Z4v3JpSikwmOAXnVsCC7p4xizrdwCb
wr72I8vrTCuL90r/oLyTtAkrqNoTXKd2vZzvf0XVnjTg7w0qiGhmYOSgwTivJ1QfRZOB5aHz/UR8
W8sQvlYDi0fWLpkNVgWdZa90UAqqE6D6yV9uRGR6KJlCPFqEre9pUW5CHwAoTnvLowtzg8Cw8HTu
L3LNZhXMteNje5TvXvgBjwBW92pZ0QBDWkE4Ud297rGIulfh36GhHJOYeg/sePvzuvCnr1n0tLfu
vL3jvIflcx7/MzxAH7+k6dKcwd+jz92foXkeMOtryenLQnhMFBCLy/ZtpSF7CPz7Cb5zC2HO6m7N
83aL2FrGcd75IBrQtIK3ZpghZWKvJInLqdu+PLg4enTdz0gWMpsb9O3Ez56Uq6hLCbCcL3SHLPHY
qm7OGySpSkmAvcDb9HBRRUNGoM0OlLxlJ1CIuuO7IHFpmWj1IIx5ZoA9YziBaQkglVQSfYa2oeI6
em2DuXtv6t6LB1uGUZF4oWgLVyXMDqR9cdYWch0XF2fkosTYeSIrIkbbAQfzToEZTUOxBw3DfE04
jUqBHIyqKFTsQ2mIzrJ7tZgnUKtr7abhlOnpS/DXHDqZrMmh+FIh/EpZQRQpUfT//aVJSufGAuQV
oAJA0Cy3QczHQrMTeZHmuyGQhaN7DUAr68Mqd+Ik65zGVfNL5rhdUI9VG7afQynRDDhxwPJMrh3K
PPW6667xNRyGlFQP5gxzMa62T5mGp2bJQt05Oq4E+4MQYd+gTnqGodMeNDYKOq1TBioz/4PsdIqa
bEUW49MkvGNN/tAJrpFKH8hnxG9HZIBDLbxyaoIM3vm1C5PjRhV9aymIBwylQ7cUEFXReyJaUdu3
ADGehAfY1r2w2gDMevWnlTim1z6y2uJcVTwOEueQ0k4XBLffo4jvvZB2Tqw2Uj8CB1UHEiDR3wj1
BJ9+CXIzTsvt4LJfHdW5JMKNPQZIzg+j4FdNrfaB7FMaTilsbULnH7/cLqf4qJ+KrtIP5Og60bGq
ToW4Z8dKBKqG2PXiDFLK/3wAHNOgkFEFilZPtCVbRhRhJs22iLKjD9YI8VAZeopg1WolWxrZdxCs
bcsvvDLgaJw5FvYYQJcxkSaDi0zxt4tURQwpcpH4+FSWn/I4P4qWhDlt3VcagGbXucgftQIAVFVK
COtvQ60C9DXRUuiRBs7Ph8rpVjFRSg+tdFiE5O2eMq+QAyhuHCRBnq0nQv/kJigbTHzwXNcVKtcC
DPgAqjAfsWyvBpo2h/ToGlDhojAzTb9B7nAD3HU9BX67We0RAH4vY6XjVcTgTOPrnw9XNc5lQ7CQ
IFjdQYlO820kW8PEwLUh3nJtpGjniDD5PqBwGzTXkEdmBm46K6svAoQ3q7hrCogaa4QRB3pY5JzJ
3TuFaZ54DruD422VxNgUWqKzWv1TPIDEoX9Aj6x+If6POXvfNaAyBkMDv57paXeAHk6oXFSQnP+p
W5LvwzW0UM5NqEuYQyWOlRVd9bJOTScc7vuk69hI2E2DKzTOCPtXp2P+C6H6TgUFoFQCQ+hLN+YS
BhQZRUtJIBvKddntE2g401GEspcg9YUBPYHlfd6hXI2+y8Dwo1o0/nGjExwpon6YVzHfFNOdSQ5N
bfJFefHpbjRGQsjIrPNXsGHkSzip61XEJTsJX/nuZvZfufW2cPJwBY5y/hwQukT1oQWlkvNB6FiH
32+j7md0Z1YpIF9pWXmse1RNNueTO0OJbwY5X3stJqTNxAwwd/rs7U7i4z6hSg534He6FJcg0Azh
TxqpXreUd9STw981HJ39DnkeJGA8yZgMVCTg/p+KU4u1z9H6GjHPD/ik77S9Aj93xE4VKXFBYoQw
L4MPWvJD/yKeaRUtDNJ8F6BZ5hpgOGnz4gBuM5t8g9jJUci+HeiWXObd/jmbC+4ZM7P0MWfdGC77
Nvl/ke0ofnIG9fzl/vq2Ol1Y/arfzhUMlmiCQfnWpU7dawYtLjBXDGNml818ElEEo2iC9km6tJih
GGpgdpGLPTiJgjni8sc9Zh62B2oRt6NuZYb2b+c52gFsV3ylj0xGWFBS5NUuA+jxFWNKkuK/+l55
WDLfU+Jbx9sBGHY0Mt2GQ5hNtJ/SE7y5TpE0adr8bN4a3y3JaPJVvMwV9QRdaXHipLK+wVBK7qPw
GDDcTJCb5vfwt07e7vbt9Ffo73w878c5G8aHY8DevYs87KzlqMlJONp6oBFByRZ9Edq6au6Vjz2s
x9vUYghFT9cX+RLrWsIiWFtKKz4c+Jc4pRyDIo+9r4lhu4wFAtqxGf+rrwNK0ELTE2ODyxjna0vd
p1mVkV59PiSHVpDMz/RiaNiODnuoT3kvvtBpevRqlNImDmskJE+3bm9KuWV74SIZ43r7nGLTZANF
icOyCgUYTfoIrlWMtPe0udvq12Bkp6PEhvXJCyNLsE1552HG2A4QNNQPnKukqkLMWDjuAuXEHxRk
srCofxl+56D+rgAyK0Jv6dVy96iogZyEoOwSCE3n76D8vSNKf88Fvoz1NDGAoi6S+QucYKgTqChB
O69RSrRJZe9bzg9xznz+Yu8pw8wU9XI3IIqE2gydnN6MD4ms6zyei0kYPKW9iGeafI5hR3z0JgEl
4Y2/zuoU8jjqtkR0L6OWW55gWWS3J0mI8FRAj7V2bAP0B7BBDRu/WvgI293rQOM6y2Nglv4AlGv/
N63mV6kmuP8JgyvIdl9HLyaKvuy9sjp1dJjVXUG+Ja7w7DYg0U6bqdM/HRD3sojrxVriZKDGewtZ
LpaUH4MgAVak2aGKAMJVzqtSJr4st+BiK9h4GJ9IArbEy2VmUp5U9GEzETkEI0BqUlWmgUokcklu
tlUdWaLgErRBS/DhTWfQHhP4G7FufY8skLRcBiFFelH2YqbXTx4K/yglzU9DJxanjYxwlZkXtXJ2
RxKtsneGhY2X3gmv49AOlU0uVejDMgVEiZEcH8HBBSQd39CPO20ZKKiq7/f8I1M0EC7DAEZlTsLx
rCIh7vw8w0S6n19CHizWberiBYG0FX3pTfu4I/ACtsWTOGW+pA+0V3D1l5i/HjW7elceaxsBIVuN
a9kj2Xq4W+f21dzDOTYlLFSOhRAxNm8Y3Pu4sqiRzHbNqFj6fcXLMKhuZQDPIWDCKGKYaMOkAZ2N
2gGC/Rk3EEOdNg3AXom+7gzRHBRmwhAk7AHbMGRaoVAsG1dWCPSVlqcdojrXObLPmvGdcZrGeaS6
4bxt5yNP1N9UGomlObkeCDKtt2C/+G26/z93WOGmt3dtIewE9+sklc04MwT/TP17XrEp5wScAMKj
3azA0GB/xtj9SIlWZDCSk0ezfCR31AGfqfXCc83/hGMxofpZ24eTqxEELFCkvrlbR8UA4T0XfFUf
K2rUNLK2cmba2nyDZvd7jkTuO+Sh6wqDKUIM/Ju/m2LMZEGXQBjdbeRdnKbxC5CLfdUT8rGBIuXE
1MjK57WSGtlb1kWTZo/48D2kd6612vjmpMEBEr9AJhLiZ1V9vbiCmc7+yEnIvAbSSp4coTVjwxqY
feucpfBrJar9vGysZ6UFAltZGNKEcJFI/ATZRU7hJE0tnJZFoWqv5IliIuvcu9ccfd5xXAQCqIt3
J8hvQNzest3G3Z2FJeMKWyLCpv5wTnfz5rZPmMA94Pjnr0H2B9F6cUpPUa6FkJeLhN1b4IYwXuhe
PZS/pOVdKEvaUbk8tv+IB3i+fBjB8ZmXHOAYWrUxr3o9th1XCtdRRSUh65HUu1hvgjgldpU5b2mE
NJuEoS3SPNF9eFH4R46AM0TBXOgBI4TGUCVxumDH7GAQRqdC+fNEVnJjtKHQqBE+BO75H9jlKCVh
VM5g3gkzlmRLsyNxPpODGZlXNLHiYNtwoD23cWi10qxNDTH5SE0yMnMZM++nV1mIq/uRld9lQw2g
tmPcaA9jsgu1pUMC4ebJBo2VztN3JfbR3ehH4wy2cmiW+CteoMTYnQONM7MAZ9Np+if4Wf/YL/PN
EDXfmmpeePaLH8B7prs/mw27tqVXMXQZcCHCWT1P44jP7WyqLbIOP3HYCuxGYU34R6d6cHHaQARH
Ff/7b7AzSlW3qmqkJ4aVUdI7rzUo1u0zGUWmsNHhDOrg+YXu8EMSyCtkPGkUQZRCE0xNIkcOXCoj
SVWRFvJT2AUu7+DQf/9OjjvZMMyu409pq0kbQYgfVMvhIprOg5QGdjTT2gDStQwgvYBvgSMKJl44
juG2md14xzC8I+l6h4o5ww/1CeMSLF60QpW+zhV9VJBJ4+8Jw3hqrNOe6Hk5zpX50Y4GDWzcpp89
mF9NrBpHiJYBgAg9JNKgvu1z67M4aNzJ2HYAg/UJkmKuNPZvXYriBM7nwEBaodSTabH32L9wDX0A
+XRgRUvxIBYk6GMJNe6Z9Kx49VY2QO7MLSvVnDQacRnkea3eom7YOiyaRCDZgnFeFoaKbWMz39k3
V3poIwkkZ6uveo/xXTxjeWnaGNQ/LnG33ZrKUAkmBYvqeWfN0AeOmlprmHkDVYKxDGp4qHJkeZbx
izQCbmNei+7qiNcgUyaunXMVlUiwHE4fmqU/Yi7TsyjRkJRSYnn6dTg7ze7F40oD20UsBLi7Xzmp
wFVa2ybdbBZzGY9TO+cPGzrrUToRwQy8ssllbeRDRGQeZTwzn5COL1NvHwaqGQo8QO6tFWOBuMZ7
PGOByhyB0cDkOBvNOLFwvsbRwNJiHUMRtNgfvVwsRMvWas5ZVlmgUJBUhjmzDfo1+N+zdC2twy0B
oPcjlFKDZoQq01zpQH6gWFq7jxPdIFMcGvfwlSmD4VwUPfb6U9YVjakiVw+9edB12/ugoyT4U3zA
AErvUzEGt8eGbVXQQx3QhNcZrwVrMK+ndTuSqrG/B6oH9hXK/kwD7XYroV+DyXziZ3wmHnMTBsVF
f5C/hIgWpn8OjIfqQCdfyIIIwdDlPurr7fJbs11KYRsz7C5OUlZgfcS0Y5T3JoL5xkyIXYs0VwtH
d490W5ST5saNPq+CzfzVwFOyCXWAhwm3S8Ojz4actAcSgfghgNQURA8F1OOOOJeqbyd8NBGIre8f
SZ7pdBLajGlE/ieyp3Tr7pTLq0vVyVQ0rKSSPVJb/+oOIPfLveeppDHOLHyQrTbi0ZLplYjV8rs4
wHo4U5HJ9bIKdrSCxP/2VFMSgI/jOmURnuUYlE9gyEK+1Exh3alrLakIGZr6b7CbjGMLblnyOY+T
v0W7LEjzv/CC8RP5VSCC79PRVHc5JuIsZ9Onvw8FK5QskBYQ2E6/wo20ZUD3f/mx94IA1+oWYmlZ
OZ/6i/iyjpWwIZg7pNDUdVCmzrFI+3JF+GRCnZ32z7LqLwUebkWwdy52KZEin5zpom8F40yuHmIm
gWtVm8qYnqagr0Wmk8Gp1i661SACR8sgJxmx+Be3+TXo3cFasCo/FVpt7NZHz7Zjjv5sdf3BQN8M
GAVw2KTnS4vOFZog3baovqNjG/uddximYWCEcLft1KTiLu9Ek9jsOhiuGbnbF5LsvaxVdxZ7SiV7
Ym8xyrmU8vt5WxHmVs+n5MF7NxEDM2s6wsnx7KUOTL8H8ZZrVzEWkTLaCyF6F+5hVaA8QkenVA+e
HDiqOPz0aHF+RNk6b4SJvXHeN7lc6VHQfcJuVV1d0xqyTzNiYBvXBKKqE8/q0e3ebKGk3cHDqoqV
vpERHihbHKY/K7uFObRkPftYQK5IDhJoUoUGoEGmt3Xpeot2lFuPdBnqCGJOCaQM8qfr4zZqt2Hr
Q31ZeDpzjiOm69Gwwg0904CknxPjerOwQd03OO24rdSMul+PxGbB1qgpz1WoKV+Qhn9Q5BHleMep
ADYEgYEyv2ocW5GmVKrzNmcucIf2URf9FvvRvXyC41fD/+300fsnTDU7ZyFltA9NIlAE6Rfraddz
hT/5t/bnvYeWCV4W0Zo7MT0dPy2biaSSzBchAp9DcR5lKJeFWYlkPRplhcERNrvv8XZuxFVDJDnu
0mDmoTPni7O2zjVnp+BImMGTFT9NkseWHp8DDJsWWzShD/6YFiJS6LpucOMjiNJbHiLPJ8Cuu1mk
uTDATULN8so2lrrkL/cvo4hoCAx6gYWv647/33wsbi7r2y5GJhc1dqpVJj4bJdAc6nGi3I7owAkf
mbT5/Zij/DHFzdw613b2IbBKo8PXvNnH3R0tnAZguBiTNhPxo4J9ueeVVIbFk8eQD+WY1hpEpf8E
95aGhMVGVVJOZpo5BBwDz37gpCHhcpEFRYaoRZVlMfm9ReDDQ1xjpoFRcxSdAX1Hrg7mUZP/zzAM
5qeruCXZcCTv+ki/VIc+kOPnH/kS7mfG653SNTtq7/Rig3jfwbViGR02Wt24xSemqBCtCDuGaL/n
hTMUCtc0lCCrjQVaUaZK3ggunUJJSDLdY87HtPMjfnklhzJw8adkuy+FPd9l9ACrigN0ZWb9AveE
hccD9IYwov9rVA+WdZoAdB1m62sN0e/ZOn8UjtqCl9jJXKWlkGbhPnuWrkU3FFj8oxNWMlhjOZ+F
MN5BRUBhawjmpAJAhYfgb7w7jaJnzSXo3yHV098HUMcT+E8sNDkjzvLYh80Nkk7SW1dsDZEiu6A7
p2AsXmWypfUEo3KicWQLNyXClDPAAp4besT4Z6S+5zpJVnNtNMKhSKKWqNJlDSL/nnQUV6EnZv6b
K5bxT6/CR+xYyBMCdPZZmeNYUQTogGMgYBigiiCuVzvYq6JHorRrt9q91/hwH+kw3RjZc3cKf9KC
hl1t1ry6HZJL+359m7JG2HIeCSsgoQu1QDyGzkGWSkDjC2/YcP/LJrAaiHYp13FZEG+t36MupnFU
2wb8dd4d9Mkm2SlMc3SA6Bbd9B21dLL4N6wyFyc+cpw+mHCh929f8j/QL2X5Nm2Swh3vktNOTlvx
2CkHsqfjTdtoqTLUkzZdAmVQtToWr4vy2/ZewULoUHo7Vp6EsUDMOdcXKSdQ+Xt9MDWMI7u9I0k3
m94KotyX45XLH7WLPJoSvS+lNmS6CJkZpVGJ6tqPzUhe4vrU6tIMk7Mqo+6EmgwsJrVj10vZ7QhS
SweS7osHkYwxIM/0Vci1s5uUMdrlmeFQJISrrBJrIFcUcWhYpjp69fPMMTriCz2nWhtP3k9n4DBk
tubNaCY+Db5aWKFm6u3D8xG1mML+9bzPiW2QnBykPuO8WbfI6gQoRQVJAX+mjYbRBVfu3A3eeo8d
KpeVlCpjZj72zp/L1i/A9+ND0Hs03hKpyk9ZOB6dvcBtxjsNagHlO8Tm1h9LUaKBNIbiAhaydJjE
dKSFHNak9IyQpzM3Yx7opZ8Sv+jajU5SBUpw34jZ2YSZZ8xhoM8KLNx2vYQtvOLPEyth4/Vs3qZc
/Lh38j+zohX/bYvoTeqNeuYNIVw1Mk/rKgGZ5aBo6ygJ3Ct7xCSvXN4hPIgw2HRskGhN9k+KFnaf
OMBsX8et9Hd0+SDOZlvyVshHLQqxW2/+M48zduvFd1wWn73mTTw+Fem4UfY2nmzs32RRDLHitfFh
opCFEluIydg+Ivq45M2ia5TJOHGdoQDh39BSsjdUp/Wb5p7ejDqrsoPXNnddK4VdsnSakFPDyfI1
EhvkyEk7ZBADWRJeWe6YG7FHMMLu8PvaOtUN5SwMUYT2sxji8O1UmXGX6MIa4vYK/LGQkFLEqIHS
4E4Gs7PsvzOD/aTAml8312Y/1tszZ4BBBhczHNT+BHnRh9Sdv+sM/3U/xPhzgLZmv7gjNuJCmX34
o4WllYinVouUzISObJktGWOQsysiKnH9s+i2o5BhCV+yA1EAXk5lOKhXsyTFmSoLrD5y0yLeZ6VS
Qot1HdUD7kJlGvbFqwgtuvZ71JfFx+l1GKhhiYOQzJsj6itlr82Zdd2EL944U30s9FgRKummfakd
wSbERBWIWscEQ9tb5S3R7ggDn/QFqk8vBmwbfZq/gt1u5ZIyfKSAgbMzz4gzEqRDat1ljv/Ockhr
3oX2EXk/6t4XDlmJtsmHbqbDmAmQAelmT5N5lBC9iPTMRv3JNvAWnqav+xAO6V1emxalPc+1CU7B
cZfS1WYrNGUlYmKvv862xkj0rS+2TGLo6TGZK8CAQAY2RpkSohqDHkH9SBn9wv2tpuvxXoOjKybf
S/vhvgRWiLvGPopOP/wUOG3fNX5sEQAsWd3HN3TXi3lOG4dNTGvpopyaGbb+oFLUbs1x442QkGKM
W11kAW+uWzLsJvfc05eVUgkYnyguB0L9NNiRZQvG+V2VoyVbwwmvmGehtbsZTwni+yrPXWcQl2h/
nRqDpcaQx9hN3k21C+GEifjKNFJ67nkMa1MM+p/bnh438BciJghbSQMcrDvn8+D1Dmxfb6UUxN2S
SjfoSEhNd/KP/G+Fu+1qgFQjF/gjJjzjl2t2HFTfjwN0Qq5EhOuReo3pkceK16n5ajTgHtczg76w
jYSuI1cSA7CgBqPYrX/jHQqqoQp/3cvy8c34nlB0Sp7pLEr15Nw+hrwZDGwrHkim5KggvkIr/tte
GZQAW5v4Tq8snXctIfcf4YHfcJ1sfSjU9Y2/XIFlqU3DKmo5ZTjsGGspurNci0C9Ocn4EvdfHSQw
rcIu58CYk8wlU0BTwDQAjYRRXDRAoEgTJWT1MUB2bFikroY6F0fdctfl0Aia43ba3hdS43KYT6uk
/CeX0nU7Gnd1WCad2yN+M4+oMfxnPMBq4pnytUAnTSawmZCAVXTlITaZQvHghM0OFuTP6G1nlEYR
orfINjyHe8yQOFDaPX4N83yKHaNFm9rVBq8kNAekmQgMAnzUKhrcbYMuutZJjq+phgUm4oisXY1m
34vwiTw77ag5Bz7Aocc7hVxaLO6FSeyyozC/3O6HzG3eyWq4bY/w1YDjDimQQe2Tng6yVexpkEoV
0jGwfPFg9+ie7S5j6WXUpZzbr4HeNcEZWeTGDhl+X17SS7s+9YEMwSZ9KeEMD7doqXCUj/BDXssD
H6ga/i4HfKAwnRyTQQ3zjL5M9dC0cJqg7AXjLE0s95w5a1Q+W3YKGHAinUzcdntlVSM1rn+m5YjF
eIUiAM3+lPvUnNUr1A9v47wGq/gOEtFZVo+j1lkRsyl9dDqPmqFvHe5zozK2vYuTkj2qJuNH0NU8
DI9vKeOG73IsOXo3nzxe1e4Z1GGblAYtmVIfneoRJCMA4CppORTEbZaZJsEIcj/NRhtoUTm/B/rE
M82mm1tFms7NBPbkr3YjQcrEflB5iDm1g5GYKoumwh/vWnSfIm2TH9stfarNoTwXfiXeDF0vzBgg
cqdQSJKKNZJDC36LZzXeQv7l4eL1MpQaNaMUNEFjCFTJy0xfZsIlQfJV+Cm12w8loMcxl+WOGkwq
zKegqwaRmf3wruOCktgAwg/G6dGKlmGpuk1HwAQcjOQO0zCKX1Z7PwCjBQz9v4nZDp9auG5mAKMR
TQ0eKxsL0kyI5gAqwHvQaX8P50MemVZkL5xzGG1aN9c9+T53DK0S/kBKWcUx0V5xRpTtMV7FNreC
EmGzTc88dec0CiconymsNUD2p83tON1NdZ5kw9Rek9RcPQPEBnyOjHijwU2BgaQsTSPfO7tSjtgJ
KNKWco9Wz+x+NJ8n5v17raXRepDzBdQmeeB4GOko+7pJ84iJpSGpLuCaweC1DEkcxxmWZ5RKKOQx
tWwHd/o20PzQFhxBW9b5BVWDfJ0Orr1CuaSF68WaYlLGM8m8moC3WY1HWvV/ZralzxCpb1TdmB2Y
n/lNaS1fNOv7Oi6GZlgvjHc3XY2cFc4tq/5h+6BdJaOerMBfijAgF5adou5v5uuunWvd50n/iIoV
VvFHv4Thy321rohRRgO+nhg/7tsp3R75PZ5czE5FNVLGi5a26IHOO8RCKUFmjDHhZi2KG9VGZdwd
HWzz8TyiYVg+vnl58/x2FrjIYcSERaeip+ViRNpm2/OWvqN9c8S/WzF1lStlD5BzifkK048Gsm7f
kvUuGqotrnlyWKc4RvaJrtwIRK+S1mipCh6UzcDts+qIK7CAm66FuIFLKWVEQJl28+OUd2aKSEcF
oq6fV86pD0Qds9y2EX+M6Cwv9UP/dpyWqjvAI8epoIT3Ykuf8OCRT2rgNq//UdiQjNmFI/aFeEic
w2G3WKO1Tyv6EsGLx2IPH3Nm/HtcymFE6ZSBD7aDh6rE/LYyxfPHiDw8DtcW7XTfAlMrJENoA5vu
+A0e7yV5TUIo5sBnU1sba+Oe+3merZU83LkgNwjD2+DxuPME8owvcgq65xgnrk+dqGMUSLti/wVq
0yQ2S4hYcsrZY7ObRLKtmCGjLPPMAzluaWT+0e7wYy3dRTLG+RQMOJAjvofe9zxZW8WXz8/qo+wi
2E5WV01/PTF4AA/A1EDHldMiHOFq5uzABdUsL2iOgnx05xYPJFNjawkEshD5gaWJoWY89bd2GA9W
P/lk9BM3aeGe/JKIxWFJVyBTBHeJrAprk2spHjsKFR4UgclCdZsyheOTXqEZHEu+zRX7S/9JluqN
YFZRtZ0jsqaJF5LXDtkxbM4Ao2lTmOakzl96bvuX6UiqR4F1ybROl98xLVufil+lRcRYWWJhu0Tj
AoCpMztaJnHyIcfs20FHV5z1vwpiQdQrOuJQHvCB7MHEnMxFHiW/cJAwK3RCSgIYurlh1pQfzklU
n8uhc/PPak9g6QxyUgJ4tDS471RlKeILF13WqTDDfr1lOwy5Y9vO+s44Tc25TQxSHz+3AsoWShx0
wejXvsIYCn+7Mp/pg3xOlcs2+DFHqDindtSj4sI4GMyw6sMVcqLdiUTkTGPvovo2TeI2chV/xDLX
v2JplueV6d60XRlOhySpRrKjC13bSWpvM3eJWTKyVDE28wWZ28aidGdwGLSv7gBKc9rTA7iLGpgw
3hTsyBwm+Z0erbAKBlwzJyNtajru3IiS8zld4NApjg9ZPdoWOlBF6Ta+7YpB4wgMaCKyXcrVvYeX
T7yEufywnFhpsQ0ekFcfR2ighw16DVirStFQGGJ6tz0HdN8wQpoYsjkNtcsBRM6e4OoqsS/Ksynk
yeOmzRO88VNVOro/mufRW+fwyRUIE8MoYNvflhwO6M7gqEG3ILgQUAp6P84oc6mxXtFX+x8wq3Hi
2hT0JIakOTzhZKvh4uWnfcFSLPl8w8zWuUmN7ab8TZoQYDTigBkAjGEsaUUQxY14hgYl0Nsghf2W
ly4ghKY7Hb7vZvf3kyF1FxnBcL/GywB06vz0Ow32kwcJ9FZG2PhJP5vp2QbCIMOTtHhkTbqCfJIJ
orv/OlT37ZaRsjrz8kl1lFWOHtwfCAewCwS1oNlb3K/WqB3sgnMFJaY70Mew3JCGeQvnlnnlStpl
bBTFlZtayaTxz+ZsXp9JtvnVWYFW1rc3rI+S0W6hb/CrWRDt+5uS9tVMR4AAEmex6JDRvJViFEAP
QLdMloshW8jmlqVrvSGbXrqHdsNkBvwMrdTlhru2WT48ZzSshl5lXgt2+1qA6NSPFE8sEpIMyZU8
dRpoh5UuTJhGuCWY00tEn2izJMyiVBF0a5kuT3NVyyuc6/b4O2h1s+32CHXniJ3u49Hq6NHEMeXJ
qN2Jxd0kD6qtk+IJxr1+AwImF+WzYa52Ro0vyustAKDWkH4VmDZvDW+3/kJx8kUY73geB8pfSuB6
cjZVsiSlRdpcKQ0349OEk1LYyzt8K6yJ5IKoXxvec6hrTgx8zrL/vZkEk8It6nWY/DU7ThuZYMAY
3WRwJDwzHX/TDA++PjlT0aLnQDMMG/E5u+mQXqFbg8aAmVf2BPfzJlyCX8PrcnvJYzCQjq4bMbgp
DA5uqX40BGEasOuFu7t3PR1KSXVwi586A4zsbInwxZVOz1WaQk16FuunrC1gVMNizq2xalNwftR+
XmItX7XbSuKrTVBJL2NOtGtXuWOW18FGJKNjTKbu5e0l/XQo93YjgnDlDH+XZGdx8pDXXp3qoKu3
W5P/3U4KUAMLLXci4U99Lw7NxnHl2xW/pfOOysjL/iMruJTCdFr/k7N2xOl5Vs+Gbr9UjCf1nzdc
u14AONouZhkDNFKfiWxzAxAYIPB+LVDc+h0W/6QHyPePOM5HPGSgKwhjUTO7Gl03aso+hVvLbl8t
HGFWiGyvCAuW8658C70p4Slfto/6e+EBvk6EIoeWx2V6t6Izc26htl2yh9tv2TdMjdUARCAyF1Na
c56eW3XZR8wOt6QOCfZTgY7a40nTKvbulNFeVR7xvKNsrAW7jIcZ4e10Gbi7WNs54nbCuEnxCwur
gN+2lDkw6PF/nEW4NxOzikv6BzAB1LuBzIfeNXxn/ITBHq+gYmVLN6fqrj83GebwzPBm/XDE+VX6
0UjAB3rIWlKai2vUlKJxZbiyUE0paKLPHUtpF8b57QiyLRQRGcXQv6oKrFQpw3R9kmn2p2GTCeEz
N3TGvsWO7ts4aYG2iZ/f83ApbGuwYYiN0J5FYKeSQZcrpIgS0fmk1850wspMiihMUgTagLUFggxK
G7qT0lOYKx0AbtivIVxcFEyHC+8x+HkRKl0sjUx/+PFP+Sp19THs7FImISulQC0Jeo5DBCfMskzz
A+5z/jviqqRaM/exmtqS5Yq8Voqzjn7NabTrm63q8RsH84UvXgVv6eK7+mg3naqFMxGwZpSgl4Lg
HvytM9sWl0SXDd1euv6a5cNvYIAcTK7jr9mX74kBhEghUffF76vO0h1PgmLp2VDC+CmfZ3Lq+Z6s
m9kDctlx4Dc2+z6tiph+fiTBfOugJ3kDCuA6NrlQmXjeYYsrANGMTBRfR24DIpG7QGBT7tZQ5Y/c
0oCzI0nCdCMTr7Ze0k4Arp9atOgHzIYC8jlbIVf9u+/bNIrgJwVqAyfElxvwf+YeDZv9GfoX0zkN
SV3A+r35mNHkeOJAN4BNjzVX2o+0XQ5u9uJO4sXqvV/68xA93C2nrtziDUDcUZ9ZnOKIf6M0Ic7A
AoTSTg+fwDiGAtUb02GuIiMN5+vMjE0x0BWek2UTlwwR8bDLnsqwRz2aeuyif31rDaDr65YONvAj
fKac1DaaDe09q2O1bvWIiI2bqkrwNw5T5wowI3zj+jIR+xMmHG7+4QF9pHOQPUJk2op34mzw6nR+
vkRbwQlL751lUyx6dZ7mxm05JcoBFRL9a0sK+mOQLXYaf3shMrFrvQBTe6djtfhqz4WugvVnA9mn
9wasKRQv6lHliKBAZ5A2QkdyDmvVKY70tqZIGo8SbKiF8O4LfP3I7aHCDH1QgJ74QxN/3kTHCTie
rdkOoUZBCqDa8HaDVOWm3fCeC6HW9tjIo/DAjwV4dU2aLuxI7kH9kHkY1CjeCXlOThfySWH51Ffw
zPQbmJKrLMkOF5ePzD9aGXENmLPmNSjQiDwMY/nA+wgPxIpCGa/SaL2OOg2e0+0pIj12lShF2qsr
7JIYU0kLrFF1q9CG11BX01NZxP/3EC0/Sjl1x4Dubgkpc4u/qcpxYHCr2/ldWnRZ3f12cBG6Wpgd
S+EnLLMi7rgCVDFOz9BBfIRvif6SegpScj9etJTmSHpkkr9LuY5GS9iQmzcpWeouqGf2yvY+2r2f
91ovfiiQMkzi7eyKTT96GtdrpQVnVI+cwkrUoxvdW0D8KHGBQcumn/zHFywfLNTartjBsY0sEEFX
rx+fCCvpi4tmkkThInRwUFpZbitYkGAVkAtpYCAgLGqLYxr/Fp1VaDojO8BOi+ZDYVs7LtAkq9Tj
FafiHh9BYeyUWAlEhjhPC85OsynVajZQiHHtK62eSED7akIOnZhLNvf9WgCbbUkdJIG1WR67nRI8
bwBMgg27DY85aqJU84XztC8klZIi7jQO5EV8xIlbL2OMRq+VLZar2h6r2hL7XDrN42DlFD1pHr87
cSOj/qD+pZokFakxwHKA54Tc7O+oYqZDTNUt4GKtAU/ty0t/yLtMKqB+lhqevMKBPxpQwqDFmyKN
RN1Ds5VCPSEKVXZbfqPf1acey/TJjMA6YBhJBGnUrucGPXi1lArESlHK6qhmxZWRi/e7Q+Vfe7y8
clmr6UuoEGSUFhLNL1aPUjVk69IAYYMPN8RO7ttT63qDzZIy0tV7okdExqRBZxMazZo4l+Vcr5BL
b3x+IFS4MkgDlBKDvgb2O4zwZ3U7vu80KaB6vVM+zDpdwGrDP/Hmcl5iNqd52UWdzHiobOroiEtQ
Gg2HOgrCpuYSMzwk8ElU1N3iPVRhfHmEX0tvxS+DqnBDPZe4poCAoVTNvHGZko52FkD1bA1eWPYp
Kq1vzP2G3PF+lC07f9uqH2BUN5yJetOUke1oSlpbd48+ICJJSwowQ+WpwyMZrca46h3gogOVVqC5
+isdYYggTULAOcYm24g2qyzVDr2W7RgPanbwFVaY0ypNOhY6lDd3AGbhIxyx45yH0i7oQ9ldKiFe
gcD49nvMEhdOzKWhroYRPPl9yV4O+aaZXcdma/wAeX27TPYQ9zo98J5bHbpFktUNZDs3ec/eUZR/
9ajctrNo1PrZ6cqnapnuY5lzIUdxTI7EiePa45NgjAsrCzYoIMNhtqazk+tvwoS+FAP2sTl6YDzY
EsW32nKVePRXxpAuxjEh9elqb1Iu7LGeF4C/klvtCgYTaPglpi+jH/jFyPnJF8Mjw+UsPgWHa7i/
DKfsvR/3JwQh/SotxDzsqC6h4hhkdFSggOXKpQMZHfp9Fh+161WTh1XtpGdADdI0TXonk3Wp3T6G
GcntGbXBZF8PBufkYT86NJzXqg2m1uYEqrxMwAl2zybtXS9FFWJxnZsX1tOmolVzG+0AR0HcZzGM
ZhIMls7v0z2MQz2btQGLJw+IN09BXG9f/OefKZ+55u53JCP+JlrkryWZf8tHo+sFPL7BtvaYJX7O
zokbQAyy7MEACLLdwIJAcOJ3K0ybmllhWqXC/pSmoq9IcOomkTwH+stywQkGXri0QWneYxTZzM60
V/3wvhpFaT2hJWHp7qu7JZAD3wXMqIf8U7r/1sjOhLoFLl1m7CKclmUmaSyr1HMb64ZTdFCNbbo9
wKh+ktt2hRrdCw1fzELNLZRdJQQtX5zxpG9l5xgLWb9JZXZ6dLGS0DuFy5Gp204KzSKfq5xaSfEG
Bo8Cp1bwjkIddTjps3iPuo6qygxWThmSM20OnXik3UXQ7E1X7ydNyAq7NGXlHygPm9f3oVwBQgZG
K+Bq4YQpu0P8Y7yxpqJJ3Z57yp51FL8PLcX7JsMricZr35s9PAE1hgYri49IgrPiVVH2CmyPE1sg
Bk7Vc5jXe/VShbIXn29zwhF32Nr+KB2lrKexqJYHxSI98lQDlty2nnyKrHAPvj5xBgKYYuNH0TYx
oJ6V7HLHDCV9mRbTG+cVHRpltprHOH2ZLw7I8IC3rbRvKYPOehYWPc1DmUzJtOhqtJ9sVLynPcaI
5IL9H4IXRjh8q71v+Ox/PLTqiiKH1fL1pULQbE4hkK/TaJ+njw0di1SZL2cbpcguv7cD5qqFoHQA
4g8Kif37tArAGLQ1XuynjPB6wzSP4SuCptlp2Pv8k644gWqqadhEVVXkq9cRv6pcfdkf45Jkjlba
JTJwSAc7J31RidOicokUSUTAlMXF31/YfMO8HsHsrnzQ8HOo2zNwEoAfsqtalY8UZNWZXTOluuqv
l6u0MXZK0MItdmDszkePnFcpa5BEgLgQ6F1Y54KzUpEd9/EVcuPLcZgdweMhuolNH7JfS4Qx5Euz
m6ty3/4lQM72PfUaIi+26iX6eIHidrattijJkeMoq2yu5MfZM0yDYQm7Q46o7+ma3Wy12J66Uh4D
O/WZX4k8TJfnI+D4biDbidqBKuNbPP36U+PGBMptCWxbDcp38aWKusU9wen3V9on8kNfXUo6uJyu
HnO/nwdxNDy2cX/XdCXYNLBqy+/mCmXT5rjTe22UACqcChMXr5S/zgCcPCZfAJUtFU5MTLQuWr5q
h7c87JVMvguxP2EbsBtTq2aM0rIRk4TBvoNsgpYcca6f3mFc+bMssXEB5b6R9wbJV4bDav8uCzwu
LTdXlBReS0kQDFjgAJLbEcnHlI1Vg1rLOwKMeMHP1QrSX0K2XwRGn8cAnLIOVXqr7ineI55iadto
ZVBdgwbB0VZ5ZhFr8M5+8W1n9jat/snKq0WUrmZCBomrU1GCDmT921J3SHPY+H4r/dMf9NjhplbZ
CcKT7h4+bJX33yshp3lXRCJSDZ/M8GLMLkKRxuBXQLIlyt40zll0anDOc+7hDfk+h8b6Wc/AfLV9
Qg7y1iQFCgllol8gXXLZOlG39Eo6mbSQKaE69pmGgS6/AE4ctUEFdrwkvhOAqU/fpTbiIQ6WOcJk
xKGEyUtTAnHcJxCMAwgBiptRKffZGu+Ei5T6wdgiaSk9IdG3m/QmlLIvKtfJ2ve+nLw+8mQiA5kd
JDQJ8jS3M/p6/Bb2kqBxD0dmWtqSKN1s+XMCpeYUnhRTKHhF3L8U9b7vIC1rzmEk2v0hmEUk9qbL
KX9/c08Ld4Uej/gROoVQkPKq+0GH5EMxljbD5QC5R9/ZxULOZF7jGvuquweLfnN+OX6kIWGYbK2R
tDUo77MCJ3V0XowBofmVHUHbxMCAV3PW5iIon3JXpYnPFR/6ytcO7FqyXEpdT0YyxGOqHqsA0G5S
gRQH5CRU8dUzLiCwHxPVXDE49my1GMM9f7LzfHwOCr9UjF8ErzAlRUAO+w7ROc/WyZ97MGBy6oxb
2guO+QeD2Wc/cM6YhkS4XUn4BLnQlAIUVjFzdAjhTqc1M+o3lTgKqDut/1UUxX7rqo6WNAkhOPue
H6gCsqEAG1c71vJExMs16IixqgxRxqRxhbASy8AChaD2KnilEeiCe8j6LqQrv0MQpYaETaKuiNQU
rZ7QR9hG2Ms+f8j+JD3QC2Mi5NMagZQ3eQlYFMn9Nq7+nFoaKYU4jx1X7EXgNmfjMaaydcq7zGm7
kYbnmyE/lHpjPUuaWQBhl15igsHrNxGdrjOMXOoLpHw6v6N3CLjON9Up7eUXYk8ISchTd3ggGM16
oNBHeMosfPb1tAoXUPCCX8P9xMEtBHpOBXstOfASF0TRMatAlo/xR0u6EBKpgDO525mmW/bszBns
RVv9PW4ZEmdazCz04Dj6FLMn9Ic46SmPVtE78hLDzX3rUpDRXysqguNpylbxsHR9Z1ZTXkFxw2Ru
MI3S2bZEo27Lg8SzmgXelTM7XN01DK9OAU4FTyYIEM0HE4QJrfQ0GD9E7WQ5vdN/XOUOQd2kp/aR
hkOBm2y2Fwkkjk7wFD/EWLbgN1GlIS2v8fn0q9XnAltoA+sOXCmBroJqb4OkA5SkWNUX/idTraN9
dLiEwJqV3OotZkCaHWVYHnHEBxH1zQYhUXPsx95/CFBDgHdwjyeTd90Atr7HRSEqGGgoSBw6Laay
tUkSaq6LvUN6LbzjANdRLCVe6r8DaWYSWxz/I+Vg1O7VN07yyqFBUrNhrdgt3lP0nN0e33DMUBFH
q77PkLQkk87f7aFCKLMGiIkUbuCqnxlCN1SSjb1ounv0VAh+zmQKDl2DozB686uS/qdv7a2hjxS9
axrBE1dju3JZladD4Wmu0788fulxgNGL64eRWDvA9LvqBQUCsiQyh58Yz9GcmaGJw92rFaWNco7J
u+8LKVU/bM+4TFvv6c4fdKgIDozH7rlcfTgSdpXnwUoYnhYe/iXc4iyEJvZ7gsV5RzMsfoaVKYPi
pNcomrTRQKeLAGMlaxtEfLuU0jQEWO4xafyUYlfGwdiHb6BqIcNwCFoeOGFH30P6Hnk9g4YBCvgR
9tW0fnCskGPAzbHGqJ1gxjhXBo2wrVfGIHMh/4WLskiWMxfAHMjzr2mT187jvaJ7RhUdDwcr4IPc
3y6gwwgtiFaG+qjfVW2zgN+ANy2tXcx3jMqYv9dsO+Hki7hpAPZ1j4M7e+LA/zudDp7iLbHpoLES
s5rVe8DGgvfZ0B1FFz5G6PMOTiwDC4V9Ptdr7quT5+GsN3vFxgoNKJpD7qsY4/4IkVpiiKv5gpUe
U6lnWxtOcH7+iKzrlgNVZxSQxUvXyElkeCZNb6/01CdUu18RfIHZmW/pvZU78dU8JPXtnrpmn2UK
tamjfmbNvpG45lJmmYm/+R4Y5XPPLyZVloKzaZe4CPeZSN0Ewpw7jYNu6nig9zVH3QSVZlybf+Hj
fCcukjxEx4BC536vXmSOVigwyqn0bIwLCj7EDYpFVuc2tzTqj4zgyHOyxjOXftAiYy0uOBe1APzI
eVxHHZ5WyFG16LX9ZZ3ofp0Lzrs81M9i9L/3QuFRTzA5SveyZ/G+YZPKx9pp5Dw5bjlO9zVTHYCI
LkxP/IFNFbswfnBx5Ga878ZNN7cltPhSyXUaKN/hcq9YSKMmT2fgrvI1g5dbGJac6MrstGeBLfHs
sxC7YD/d4IjbnlnxFPmOaq8X2Ss01+L4cLUT6ZhurCzA7Dgcf8GL8wvAY3xGI3bxqQklNZXvA7b3
uS8AixwTFQ7gT0zWddqRLZj1mQ3Jc4o4u2t9SijuY+QMG5hMk6BzHBr54ZB3SLTSA1rKxJXZSgKn
T2N4pV/MOpCSBqjwKJy28Yt9y/upRq1gV+1OYwydz3Cbb3mkUBlXVbPNF2LqkyqdiT6ZoA5XNaHX
bjJ9FYhFrhyCA29Z3AVpLNfIKAG+Y7YkAKuiy/pKVP2qHqf+GsweMVUyB+lqToKLFky4TchMr0N3
peSt2hhUfhKhKISk4WBMa/9EdnPA2vkcGiNs60lk6JchQyPoeIAc8SXZ52+zVQeA7rIsMGbVK1cq
gH2/7sCumlx4GF5hTm53uSuzeNncL9wXuSydagT4Nw5IwVhxmpmVOVtZPVCBBCQ8qwl+Id1sa4rN
kHhjm/NPaGbtUTdm3lMEyyP4sHdcSJhwOcfrUoPYQSLWPf7YC8xCHsdbd9PwbQddZOvedQ0IwZdS
qMRlItxAhqczEZKI7LsJo13t8RostcA2odmbOYc1Vyk7D9Vk/F3+J8lS9/ZkSmZ/PLMXVnrSGzGt
AuRP6AnaUTg2BeMI7y5QioZ0K5xU1dx1zhDE1Hurzl7IkQVqWqeteyDvxqkpf7IsUPAAxAlOK4nA
x3/AX9rGbIdKeTSc9ckjGBES0cmEO3Kuqck99G4FWfTCBPb+wR046YBXPs4fLnH8NPDNdNV5ZYLW
cU2iSwuPpe+M5fHB4Xzg/M4/+ZsaqxHA5iMhib9NpJZW0TMPpkXyZMtQJn+suk5luDWKwg/zvCr4
TeuLWU1f+oarxo9C+eM65pkUIhVjDxVzpH3qLKxVv0eb0wUdog7qNUEb4Fs04AnRot7gB0FdatsO
W4+VLZPK4MdAszF+NRCPvYmOkxJmBM90JrMjiG3a4Ael1/0Ho8YbSch6Nf0OzDgp4hpcqPmIuBqp
Ml+hWJuttoye51CR56NIjlleeBrltmd3KqRoJQyTxCZm+UomgvZXCJYnr5yvMYDso8VR9QJRSa+R
M9AxZnhTa5DHLE8w2IZVcFTAzB1B812X2sOlAOtluY3HZdlJLP4JfCf8y8bGdmdV3e3hmaCZ+A/g
MKlFtlefptGD921VBgfkKb9K7jEwQsjmgcOhQkVwsGaJdDxh/a9KFkGrEdiYvGWOi6IX78tQUk+n
4gcfzt9KzJ7o7725xxoElvY1tdgGAL6+NQ340fmdnwNE4juanMD+Y3uPQtnP/YVD8MCqDxCILS3t
3YiqLSHzPEda2umg2QtpoSq29iB4IFIbBBgIKT73UITNuILdlLnUwLq6eZMZdFP+Es500tdOCjar
0pQmIdyFw/j+H5jysiNG0fwbi7VSYb/rff745/XXsT33SlE8QjNdUOi+uU8jKLG9HrOstgAGdr4w
PrAo7NMCyzaktjOZHb/urjJW9RKzQJzj6mlqjd5zfDezOVSdjBqUsnnvYKNnKMlvRd/tcSi8roe/
V9ZOI7Kdy2dycPaffQsMf98aeuP3oFR1ecLUbtFSEMUDs47JJjG0lkABbdu11YX5zhHUPyffsR+J
myCE+lxTr+eNc+ayd5x+bOLasHYNc4QZo1dbM1wj8s0ZSuBtJOqgiWk49OSwN98ZiitZojaCX5tC
eheq1Z2QOIkrTkE37aNPa3hG1lEdwB9c0vYTdnGIVvnBdZYGOafzrCRv01JVPX54KQ1omo//qh/i
fSTz31eFUOKg219Nie9ePMsTLKzHWiAArJ/LvXxfbQ0JYtBiLNkkxv7/pXP3NaOmzvvK+cKs26TA
mnuGt8BabAJxKOaF2NVyzsqoxZO5FPpK20iNNHHLy9EwtfdYkt+I8l3D89WOQ4M5umypMaoIACAQ
umbYCzPN+YTQe7VH/tJECogpWNB6JrdIGmtEHsi9kgAfzxOh9aDvmo+vALbFzdd6w7M50BfBsheZ
cXvZh1Um6Ux8kk++6exS+BrN8l2RAFjyeuxDj9hP+1FRdIRVhxvuMk36UXOxdywvmYrRguk7Eh1q
JNg3p9r5/Kkw0IhitvFv4Gu4xfdcfERT3IzXzTWkIL95qGT7nRYLH61q6j6bv75oAyA9PwkWwdkw
Wi4Ok8p6yNp4F6plZKi03eZxakNbxM/KKWtSMESQn6TuSkE2Ag67HGAI07AjC7matiCdzMuTt8Af
gNCMVvEfbwIK17JklgWFEXsetnuinROGHqXbeN93wQZScbmT4QU7/n1Njub6Y9gd1bHk0aUjgm3k
EqueAfq1fEYjRmsqzSwqyF9/79d9sQZYrGDBwwf148hyOZsd9+IHTsP2I1zKeTj2A4inF8c/7bZa
5IQ/DT5XSsvawRzGMSEl1BotuAJmo+x49sMziC52USzwEq06bVjTT/XC44TbfUexQe7sjP7+SW6b
2Wlrp1FhGB0Fow1weRHvz//1cyxwz5KKpbSJPKQwvuEMEVflxcO3S9QVJKnkdWah1H6MgaCa4PTN
HWBS4NjSxr9n7J844LPyvN61umI87bVDIAznLzheBQkqmaSn1Pl5dRovzMKPeXxt6oxcCiBlIcdM
MuZQB3TvBF+C/jSs4CAt8FgBJ0/gZrOfCNbg0mUK+6rfHfZj0Nn1y/wi3IoL1DowxFKtzg6bNrdd
wJB8hyAOw5WLStaGI5KL6ZJihS0Bs+RFnIUtLfFvl7zR8suZ8mCAgFVF7lZ02ADMdYbuAA4RTkoO
qbeyKr6AjYte5kv9EjTiLXHDzo5qOgpCupwGbCYRGeIwfIlj2d2kRpF4FvPqP3qicTkX5YU5jVvW
VvRIQQvYnG9n/Mj7hXncRtE/mQoiGZjaNXYpIDaOM0HIHDURC5p6yds6zdtNZhmKXlIrqwmN+CnE
62LPmR0nmRnuqTNhjaiRrRrOqpb7ogkZL9nvrNHEdxmFEv5IjXxTFb6lr5P9htNNM3ghq+36uy+t
hq4WyDTrrWJXL1uyNywnsglxQBiVr9lPO0t2pDsxFj9GMAi4lbGuFkfm12neI0UwEMe7aJTZQPAj
xGbF+GnUK/jE7hkSNMFfAZP/HbVoInHEzWS7oMXtrFCVkjl3GVw4CrTke2FJHzuIjO5QfYoCOGvj
FYZi8KFQu9hoTIMLvvHr+zkOj2yHLLki2z5M7UbMe6pRXAxOPQ8UjNKOCl/QoCZAhroihMKOT+XA
I3mn0m5Es9UIolvsdQ/Sk3dePu5OH/HNeI6lVoRLoFgCUFT587fhC2ZTXm8miWU6u0WNLLvmBaFC
1KmqRtmvq4NUphTMS75FRZLNIMLo0mKxYgXMMOU5NL7QdqWf/fJXKx2o8HCQJUQvEoZDVnlyyfRg
6p6D9aAMI7+6wUwyNjMBKZj7wsUsIraSaK/sOGfQ+rZCwCO02Ic7ydtdUBfXzWc0kHjmcvvuvpIL
KtVGeq98iwCVjHlDc/0FNl2OeyFj7mczwWRb607ASOXnoR2uvSnyGnWMuzazCETLE/uD8U9f7tbb
y1FcbT5nCcpQPpwQv9TJAVrVNpMXqzjzWpjy9wm6b4TtMwZiW0CfNANUNYz97ushGd21tI2Qrpuf
2CW74OWoRwNoUTBVVMdVCdkxYw4LGYx8inUlFdWpSHXYRjAC+leNB/PEZbJ0Ced/RvzpWQsI2447
lAaZgzNd4zRBe3Yz1827o3o41en7CT4FkFLi3PrNddYL27l8TEZb0+sehK8hBoAbjlRN702+SbYg
eI81k7Oxbav/5M5cI6DPXXpN6QLSM1pwjTbarctwfR7q/hLaMsvI5CF33t05ShFP33DfA6dyC1Jd
enLOq3GCk6mbPuE8ZBk9cIbp675jWKggYHf2YxZf8QEy9jk1ii5+GKM6o3qNnXs3tw+jHaDfMSU7
9xkFL7GdfGk8XWRvVl1PL0dxga8pJBGZKZw03Kr4TGoVIqJl6VoI+0EcdDEM2WanvAQw8/GUayvo
LYeKbYwhaoUgxxcp2Jb0UBz5yJdWJqO5dsWewj9NlJq4jYSJ4wnrj82MOO97HtmciPX287t5Vzy4
YUoGClywTsYrWpLD616c8+2fOMFzdqFWw9Uvat1ggEP0tb8CB1c5IDgVvSsXgPf+VieCsCREnziP
YZbkHkULg8f3JDa66Z55slT1yTSH7Ioh0Qg7Qt1qnSWo+hz0OlalUaANYS3XSfMVWqdHSb/5cFID
voCdk7EL9qsGPLNpZz2oQL7i+XnH1R4cZFjN3HVplp0ki/b7rOQgiRvHvcHYAo821aExgE8tMFR7
Pmh4b2Giu24SXsexLnDiypQLGcUjHOW/k+Udk02WOiAbrsN02xnpUAIL+Z1cMlse+XfUImWGIdcD
QGsQxeoBjbeoxJejCkfdVTz1MYHIGrkdb1xfhShG+LtZTM9uOLYZ0g0edcHJRkEhN7Ac+6LP5ZF6
RJUD/GVfXtq8YKG2fQRAML3bsvrAXnK0uNTl0nad6g6GgGffALvpAGnZSTyjvPP/2Nm+P568/800
EriSB6aqrPTJRo9xlmTh4QbZZlHoc+nb2AKj6zzFPb7wwA/uXxs3hUPpLL8Nm0S+dX7XdFLWNtfd
3MU9tsr7jVWNDfE8LYHDTtmyCm2mm/h22NQSpyioieR6aaN97bK0zF9ZmXLHbAmF9nJkvpFJyPl7
N7AuvrzICrWAONHfDbqJMOe26fxn9chZQ7JyH3HxXHHaEgtiSLqMDAm+ZBARvVTUq8QtDRFgbsMn
Ik+kKLuNz6QFWr/O6MsOFcpOYLDkwTZBtqLM8pYfNVTpmyi/Lp9AhRMCIoZo6CkJUgS2KvZHXZvd
yjbO1y0y65UhWbHWTX0dDcv70gLL9vUjvUncNBbLZJvGXlAQsC29mghssm9UxWjyTRnEE1K7OFmj
IWCjuFxbVyzCmcQ0l+P5+HS3nA5asZpUyzONxBhRXXC5vaT6/Ws3ioXkJgg8C9cK64RfKhMC6KVn
sWYoY2Mi/U8dYPwIyEFRr3PXK4KeDqBA/l0Pcf4AVPsljcNX9VppwpL6xqSsq/DsUhnHGcfff/N6
b2QKfJmBYoRGSCwvbi5vrI/c9VsjjNZq3jODaJaNKfUoPnCqeJLD6q4r4zgk+uguvDLmyUUZ7aS3
v4s5zJYknaUXCSs/HDAukfdPAiPGXRjwuA2XoeUvOFGbi++Gn9oS9FCA8mOnFn8qr6N1D16DJASX
KlR132vUm/u5SNVUD0+Ur4rEFzOGVPSIXIOmzkFaqhc7LjSSLXqX5cHC6wzbHUZzX9ANaZgFUxjy
5qCnXX0tGv6PnRIXr69jG9KIZ3L9xfhuw7R2weUsAd/1mvwy95W3wyWoWxh8C1TzX16DvPZC1JSf
8sgW2SCPeQcZBR4GmxkfrS2axeQLXdf4oUKPWISZdMGgdquf5LimZ5Mooa/VNp1LDMEdHmHcH1L1
TlPqmwDRfD8nbPLFGZaGA1iZ4K7E9xR+rPvNgK/Y4JTpb965pYKh+EMHEipW0CVGgd/DtSx8V50E
9NvquqiwFBUjJJq9aNR2JNkdbRMJO27Kyw1nMBrHnJgrAWvBln6Bwh94zOa1hlVTk8Yo3puqozR1
BHvDR5gUmKGVzXzSZFIXV0IqABdhs3kp3bXYuJHH/ufW2EOAiZeyZ87o/5uleCmhPt4SS296Bz+R
QsQ7V80nbtyXbRJhFxXhmh5k6GYTzUhLkpZSUtHQx/u6Dich88Ucc4S6jQPLVyzn9bgM9lMRL9FC
zTXpYKG9Cyd3WOfU+FAF2cX7L5nENGq9bZEfL15y/UuatUk0bl3oj47esdn4cJBNyXWsN6zHqUlg
DcriTgEmWmFy/JNNA3IJKO1Orrqs6y0F1fvh+UnuRR37WtCQwo9Fn4MPWKxaAoXDWlWZlTVckKLH
Fn5ErdRM6vRF1D1UWzjnh2xMGHfaJqbhTWEkBymHX2QXeqmWB8Cc+3Zj3gtqzdFJhye5hLW6iP/t
sTh53LE5H/Vwd4JvCPFVV5mbYUhWhDxmMiRrnqyw6yNwpuukLeZ6fuHsWpIABYURBMjPJI0jgrIQ
3V4mdUl8VlrvORLww+4pjPBm04E1M3CG5qjzyNlI8gyb/pJFOjt/tqLtveRxIckW2Dc6WRYx7NJn
alSI7D8TP7lmsqjir5pVFtyN0uzXut3b54rC0j33P9I7RM/kJ9htqGwPypaixilxF1e0K62ty5m3
YmC1dqU6glPiEnB4tSlw6h2PCZ6LqzSGislMjXR5uBNIO7Sp8rF8P/sIRI28XQnkYfnYN3eICE/v
LicgayHB8XbJKCvKvbn0mxeOzHh6638fwW8gK3P11kI54dTIMVH8fyoLebnUVU06ztjcWomFsf89
rFPtzXcq6nXF6Zfr8aWmg2L+Funa3sw0x1Gek0+cC68d1V962LRe3JSlEAOvmvy1paE7a/cxKChX
jr8KSJyo8Wt0v8LFnGXseriFkylPK4sMCNL6SGjx1bL8Heijm3sqXEWCpzINvnP9P32J2/zVSnBQ
kX8vNOq5q94QFvdxpESFC0NJeKmH79GbG/1oUSDNmSPDG1WUjdaatrpgowphBM/Hx3+1YIrfB0PC
svF5Pztc99BnuOnnL3dItx/fOWHWhKW4S7Veg7jX3u5CpXEUvTkMOFjn7j/uZ71l61u+6uhkiVzH
YhvU/rZFb+5D80EPeZq4QYt4WKLuHmEUn0v/WL2TIZxyaSskUNXGg+3YtaUVfFru9DgHentcp5Q2
eIj+SyVayq1cR5CcXM6zKr+0XyEGyJGgTSA55oVRJikDOPeIBsiMNwXlJhD4fvY6clowpHzYVaPY
f7c9camsVYPdiR+aGLtWmiQb7BFPgKltBydZ7by6+NUWoIneJXvhe9WgsKDHXBf9bUcf9irOPv3f
PHSHiy4t3u6OhXlBDQjSh58rJNANqmxDzNx7WXI20AUaEa63wm1ynHgC6jUDUmMYA22bWMSuXSBE
H3eRxImlBbBF2S0odgaJXfMoF4bp9WIUNuZ4WLf9v1jj7jCHqXIbisezYg9bdnweoCt4wzEW55eZ
23gkkMOZN2jAouwfT5hi0+QV/fevjZ4MOngPskWW8jS5hDbyv6uoPLbw5eY6tWAeREMVMwKXJFh+
xfxX89LPZ5UqkgPDZ4gevl36Kb8DWcdpSe6px0bthHQWmNX/n/DHeDHW3dkuC0OM2YYYG8W3Awqo
7nbAOxd+8flCaVPENEUg0tpRrkLjpgK0TYYGOR2VT43S9Ti9FwU8HirH+C5tY3+zoVFgx010jJyP
9+w+PCLoV+YuK3g+WltxYH4j+LyskEK4Wupv9kb8dsGdNtApZ/w0BEi40PGErY1l3v+8JiKcTsus
rkVZyysB9bBkAEex6ENrgL3PY8hP1c5iuGKjQHywQf5SxQcCrRis5PFBwn/yhRJVxbdKjKtXqhY8
mZYOsTmpk3n87Xg4xEiPUWl6HG3pZNwEjjcEaM6+HN8ttxQyNZwPatWwVAFB9GCLYB/nOV+PGjql
oBVnio7PVNjuYLlV+Is138Et6heRhJqObMYriWaCPJzO4gScw5wpB6TzbWMptO4WvWJ3sTa9fwWs
CvYY+7cLMDiNN1iHrzsmFS/m6OgzV3Jvgd4jH+G9kmTwNA/tw7xFNIK0+DYeWVMZRWwFgIc+E9PL
cZjfACInih8c+IBU3rXfdpNWL0QJvJyC5GXYWo8bao76/k0INLS2gChUYt4dOsd6VZzbekSOah2S
l9eQQUa/VU7iSyPaD+iL4vh03ChtGWwsHvZefDLH/t5B6gYddYbjPsM8v7OFOy2zGkOROeLXB1dL
cfCsz+e8/1D6kfJGMNwfG8n4x/h4abg9CYSl47tp/MB14bR4WENlVlFuPigfXXI6wuEN3QQbir5P
2aOP42zeCD4GSUQap3ZfICxh2Ke3xKugb8+wtBrToQPObtk6ZnSKnB+p4wsohnWMXZzV70E8DZWj
gGITe6Uzn5TlWae4BLoHhmSu1XVh5GxPePNY/qitjyeIXl/GD74l2ojXgHq2pjT5QUVmgsz+Wwtz
GLRsBWGmujTv+tYGIq4mfddZbGj0fFtN2Ci7O4dxPnYdKMgsrAJdO1aGuV2OKfj8wVmRq1bQDua1
sMG5Aaxeeu8mK8L4NEqoLcYMcdEYLwTtQZZo3rBKp0W1lJRR7BjVLpmk3urL4I29e7ijFAd3zmyA
k3i0kVLwQ9fZqZqouWsta7QCnCvOsntwfhqv9wlCevXd7dP1WJJdvEzfla5xqO7K+rGWIZJs6Z7F
DPKWoETfSXbsCluaSZ2oHo8BHYaPYdo9L8ToKv6Odeu7ZpCHc8zGu1+I2NvXeO6lwhkCDFFoNQoC
eoTZr2nMhy9hetcCNruI/kTpuEzFMaXqWCfMxr81w9wcsODAJ8wYNo6zaXOhYKGcwz90d1MsoqJ+
PHHSF4wuRmCGpgtiWC8aPhJf+KAXb+Kx5zaYMT8musL0+44hE/LteAE+ZyFmLoWu/XOzCjx650C/
zhkgpncIxnldnYto45+8gIoK0nIkgcNzpft5fauSJ9ha4OHHANcDhYXk0gQ911V51UrWeXlgP2nq
vNUtbwl5txxCc++fE5prnoRHTVwQorCX6i6QvwOqzOMoaJdtcSKiQQdaxTfqxNb49Gw01htYVRv4
hPGt7Uc3LK/Q9coXbsfpwLPcjI11Y5ABrxLV65PPhc3GEboOQKmGs9ipduoF8uBegJ5khTg324ba
Kx5MD5iMVGUf1KDO9kygACoC1Z8jXyaufXosK5aakpWAcrCacfge6vdKswj9d2/bX/RGSiI5tumq
MLRjxER3Gp51wyI9dJbDlJV5tu3yiWFupGY+5pdDoUQs9iZ8Ge8odI6EtmOBEEVBThPdPWbV1zVJ
GIsMT5uKcc4J6/2jsEeKMajrNgLjmRlJkT9zqhzYMVvbg9/EKa+mMmB9YjWx1n67xzyJrQUi88kH
Cqx6kp9plDwiCeBi8bhrgHD/vjcl0ksReJRncFJ29oqxJVqly1OBLJ34/4xmQOI2fqFVYhDuPHrk
FZk0hUuX9lyTQ7SUTik3qEID4hLPMNaj/qKGDe/N9dwQEKc4ZR3HRr9dwB6271pVgooq9+Zr3W8U
U1/RkyT7YJQ+fFUP3upsGpiD9Ab1ZFH2i9euSHa7/WOGRitPWs/oVSlXm1seq7dI5CW6milrsM74
Z2MkMLlB0qlF/GRR24hLu9UgfouxExKWHDR5VqR6iaKCOf87bOmku32pY2JFnsUjjy4WYF10dYhS
JWg51bziYKR+AG1WwKcDokc8i0PJkL0dhCrTpc87gf7CVTopFhXcbQ4aBJYBNPlK6RfvyI6A+TiE
K3FN3adOc5YF+ReTzuclJKJChgMXFINFZBCGk1rjFs+fV17X1aYiQSnPJbXbeQEoSokqthPNzxBB
VHn/WYl6LxcBVRX/J8npkY6foPAnyDiIOv+zHfibGC2ala+j9+FGcM8zp27dRsgdB1k9vM2kNr7N
9wNzpWf/4Pb3GH0h5pMN6KQvkVsxI5gz2NV8CP5TyJ/VCrd/1vqIkq2EKu/zuVKeG9HOoF56H5Fj
CuGqA+MC7B0CsyW5tbjDwS7Ebn4lcvW1CSb/afrDEb2T/+gewtE6JD0l2Dje7LlYT1MGuL3Y9Lb/
ev+U2vFZMM/R7KcLxOGb2oP28x+20OhXi8Izczkdoj2ABV83Xeibbj3E5550Gf3VPWf69OUTl9K3
TAUQDg6C0/aS/WuPDBINxoGby7EtEVzqq9BqSJ3laD7AzngWDL1WVZn2htwRCUsTTUVFQfH0Wt9f
VL5cqzKZdXITL/T/ck9utWTwhSkGQNsaJVnW4WK/MFJkW4OZxJaYMZGpD+dYiPRALooUlD4Efw5u
hrcTUiWfpVQ2Yk0dQ2pJLV0xMR76HZyhOqTEO+LcnhaDiAmzv/v8TdIroQPnqOJBUyaVKWqOBdf6
PX8954hyXLXVwilYONjyvjjtBUZF6wFE/g6ViOw94xJTUhN8z79eYYhNXypsLvNhzzXWh0/YzH9l
kLDwGTlrOjIedCx2vmEisAbaaBTm2Ww7WcZq/f97YtgkxMkifdPBMpXvC9sn1tYsR4bMTvXnhFf8
3ARTmfZXrcIZdhzrMj0GY4y4DAMnNFdlcCZtogjY/ZJoeWaBmFXb11NWPHaTbrhrr9BguoGgndd9
G1/8l+4GWk1DupJOSk11c/Rdb5BonJFi+8oPmOoPDFogvHlMlnBh9p23CzrARiG/mIbWqHHCkIQT
a1HlT2QMGNkAgrHSEKWcrL7ajGQcQro7Rcz2d6GHYjZqbE6QwBtpIWWBbXkbEcoC16Dh7mYm4EO/
n+HDrlht2RbalIFcZk8r7bvhBv69jTHAPEcR5Oe+fMLpU/oRstDooJDMuWUMgOUOSVpQKPxfb9aV
2Rrn4Zn+pmPtJ+7Q/vZdnRWuETrt3CsfUxFpIz+xdkJSOd/vqNzC2FhTNIHg8fhUtbw/MuYKFcXr
YE8fipnuUmIagQprJGjs90j+9WjHOoVpLsKBvcIDjgdzqJGjxZXkLRJtqepT4AYy35z5P1F5JKlj
9vk7wVkTAlxnIvWfI18uXGXsQlrW1HqiI0MTHzmzcmzC8cjvAU53UOO4WBj3aYSa+Eg61YTwsKOF
F9JKfofYo1Z7yH+zxImdVXJf+P2Workx3mCZQ6FRI9vrSAGXXHzmJlP1oQFMkQu1gvg7tPGvSBRe
PZnjq15+m58Usw5ruX/y/epwJPLXrIRmUX2YUzm1XKryhH/A2kdrf4lgyIQC9In6puW+LXPSsf/u
kFXGr4PKXs4ZsJUEL31mSYsRIXz9MiWT/vENhTVW6V+Mm5+VovimetfsCP+qYxSuevyhYAgZWPY5
6PXU6b3MJ09Zp3ReMJzgLZNHygmg1kg28cerFd8y779tMo0U4O6ab426L0nzYFHn4GPQ03CcmKQM
gwN/mWlHDqAWI4OeECxvDckYcfHsZpFS+tBc2019ZrWUwb/O4SDWRc1rgwWkJ8KYK5AQxYiSq8R9
YlKpHL6PQ9vEU/bZ2EToqQc2dcLjPZEHR4K4dY2ZW3sEUaSztI2ElH+Wg4hBtKK3KuvOBoy/WW0w
yWYpcz7l4tDcr9neEhi6nhclJf/3snwgVHa8bWjVHqBwbNhKpNRHANjwWlypGG/0slTJAoU6Itg+
Pg1j/7QHurDm2JfnVmTiOkK8TvFHKTMI5s5Z2lKlWpR2mFaAZzffJYFZujakhihb2A2W52GI5+Kj
FNvC1OolNyPfCXeuSFXBcOngbflavkS6SI9Y/h7Pn5M5ZlMeiNVtEeZZjkmRegUT3wZv9wSJC+Lz
J/bUS5qN2/APJpjiC4dDPV3pnjG3X/9H4yj4hqzPEOb2cWPGwcCfRHIrLcuZFK3HMreKJjuQA6x1
fTNKy0dHurV9+8Hcy1fwyqFvWAsuuhyyZgnI+yya6YxMrqj2x4Dh0kF2KDcD3cc04TDIa/mEaara
DhJiyVXRRoKbQlUPNrz+9LBvFI9Y5XYZzxwewPPxGx1hxl6fVaTVB2UjqcZdIzZAxvMU7kCyc12i
qeewawX6x03GYAM1xXmKAxy/3ibyqhP2NyhvZQQAHjQ5wqmcGULTy5wqjpEMKDEkqPA77Ek4UEXA
wylAEmSaWiWoN8bzBdcbJYfV87bKKZyu/nS1dsGln/CD0UFvd6+/l/Akx3SihlerWzFnvNcwaA9f
NPZt3T9ntC3t150qktea3HAJxc60S1LAckOlbfrqzdViwihnGXzxUccyMNDEsj6LEk4y3Tf0E5lH
OebVA9mRV/3wETR/ij16zP72ZNLoQyX1X/IwtMUUnOr5H1cT5ulqDbi6MrtrlZ4OaY7pEjP6YxXe
4arEKstZ7fDzSL30bKYPwXlLWqeLEdgFIosMpMyRScALnJR/8o+AaN3mwrvnvar++3IGJs98Hons
CfKRaAd0AO2P0zYl2a+tz0MzwTYjX3PT8d6H5Vr1gRPF2wJ9B/dLmnV18M6+vkcImQjrYyeHO22M
A/bD7DfgsIb6ztTr8TsoZ8QlkQPQ2q+NfsxGAt/6JPoAJNFCSMVX7UoEYQUKmuNI3pn9Lx9XDfdC
FfKY8SohyzRAygX83pjuWlxFBwrMC6aYnvh2wgEguN5R9x846ivLF0PVSKmO/ooTn2ERVcB6PgKC
2jUr0Q2B3Cs/LFF+truLv2an45a0LsfvNnKO7SLEXqzhKmSYLP8AnPTZjbFq2pt7/Sy8lI79eWM0
3MGM0d5LwWyeckS9EccC4qRyXvVLNo6St2rirzUECuNRhtvD1/Ib3kncwaKdDEQyLxndy0nv0JuW
FbwWdSntZvX3vEEuHDH7r5yltrSLTTqfwRBsLlatgHbHrtO6NcVdbI9RMor75X4kWFDohTn/tu4k
rRz0zZIuubWVJCk5k2BbXY73LUZQWLYIah9nlwmFQ2YmjVSALr5IP5aZ5N6S86FvXlvQVBkq9qzY
41PGMCnSYqVEWWP0t9KvI8V3s1A4rAKWyyQjs7/52wtvY5P6XOJlqp5I8kSo7m3HmN/AlEkSv3UR
2SJIvlMLECQEYIwBm5Td/mJuqtgWAOs8CPYXjakXxb/ks2G6DqWpBxLLTqHF/mG4OfVj/IiOwa+z
g1dPSmkITQhBEAObeab+lwMKDWoNDKluAhVT7qC8dm2SMuyBnqQekQelrAt3m2EqcRd6JRsiM0LD
j6IDgPQj2Z1Bf+UWHv1nwgSgfvGBa2rdc0qSaFdcZYWhqO0WMskq5CkI7u6Vby0wGx6uYyLSZoXo
HOX2awsGdx9/k91/zwMEg5xsPqMpGYMIusmA+P2GsgfwMdLdah+y13YNLLIAIgCRQEq0MrPcMe/H
AZJu7iMu/TM6kxS/LcALsEY/ulkQaI8QSAhB4abdxrwl2ygNbJFEjldpRGGRVcYOZU/ZtgrVl9zz
egd+uOmMy8ZUTqK/da2doMU6zDYLBemCNlXMq55RMLlLlow7kwLlxvRtYE8Rm5xRyjlBJPmFf2VV
0EY9lYS9C8YAtgBWoNyOdwh8b5CYhACQqFXLvH+mjc1J81RkHWBQz45aAYX1Fk8uxqK0gzjchuto
EQ+9Bds8cTQBDciDspqddX8SWGB6P95kVdDk0jjqgejR0zomgsK/Px7HUEfuvrr1tbQm0vJkSPwS
qQJrVWL+s/v5ARbHGPL5GWcEGY36/yPx+BJ8iAMNWSLS3gnXQH5pejTgwo4i0SnJcw7o5JhgQApB
mfzzqgp5CMTnhNvqA4jnFtXoxleC/NkfLKJN/MtMkXGHB9086yi7PfTplZvCrYpGPNu7f8iO1idk
zrdYrnojbvjWbd9F8BDptYKrp4souqzVcj8udhxz19QdlPBPyrSNHKGY3rnst0rt2Tosn6GeCj4D
v1nmX7fJ6FtuJvmrWCoMtSQAmIOAlaJMdc8ZJynlJVK4qtTu56H3Of8zbp//vpYCQ9o4Q8OZQlhf
kvoQ89Jq9ngv8f6lfzt/J9ipPjuiFljiGIObll3pseRLhjkSkTus7A1Zn6YTasS/TVY57vrUcCi4
8ELRLtz8BFsWid5aKWmF1smnB8gzJG0OYFsx6MLQsvx8npiDlQGvRfKZZsAEuyc/dWu71xJi0Fxb
NmF/FJrD6Aec6gvtPkro2IseYAhxsUTTzpmarfNl1rft6W8urLE2fYlrQWXbrO2D4qS6kK7w4Zre
nXBfgXjlhfphs0ms/tsvkSC1VWY0tfnrBq1t2TSpLhUIIrKolYpFecjEHLzC4NAejXYceUsKztT9
FyCdux5fe2AbUFEXaOuAeR1Nj/dvYoDBPwbgGD1l/qDNHb70fM+fo6Y2O6tDj4hNlMXMtDZKS3OY
1MfA2qEX5DlWEIuKiPfY5xYBItUU9Rs31hnhDAYRVuXjdZHnPRKZZWfa5MgG+qTe/FTCGwJxlxcT
A1Z4d9ciBTipy99acwjGHv7ghbLWIzFn6llyN3AMmq9LQax2ilbaatMpYPPUq6F8WSmLH3x+xOMl
02xLdOYX4FUJX2C5wyhe4nTihmvLLmcfbanP55OfzqTXWxJAWNxNB5RhakfjYknARc7zEEEHAsiz
F4daKGexCsQJD8cwilDkhYmlDjhCAtvY+FFqSnS+perjoHSkNxk/wvlqOfcRlxhNIArzWakutrbs
UwdWuETRMwt0VsdhGUcOH3aH44ilnBelqV3Ecx4PLopoVwPw8E/7BtwxT/QNOkQUwj5JDnyXnlPZ
+iuO7hg0d67oXPGmvb7Ktjd3DCLQ74NN98c/NtgaPWjkrE7sgT9EnuFuzaDu/6AEOYxDMc3YJRZZ
67CdY97yOSA5tB2GSeUW7zOZs07PzAQbfBioYPCrYq7jFWK/xFBFHXO/ORDFo7RMIX5LzmWgYE6X
7bUp3pOTib78oCVPdsykNohLvAsZD8LTfRHB+8Zq/bpwk6wicXc+l86r6HaXIsoyTjZzXQI6xZ1y
2A4WV5Ku5wm3rhJpIt2wc0Nctv9dUEH0Ld2odeyvfD4c6mrAFpFxC0TYuR/1XnhUBjLRGTL703Y3
Of3kCqMCWsfuj8EehSbXLcRF9bzagiWVYH1CvV09Duh/9iBXSzOGSD7DXBqNynRAtAUTltkpuir3
5fQR2sAaUAgurW/E1wUYtfB6IG0Su3IqdYwWTulm/NESS4XT1atrp7moTVqv82M5JDLyRH6TRu+B
hXqVWHSj40oYIdMYvaX59iiNRGQJ8G3IzCVSQ20bGlhgN6wru+zauCTeWBM2dc7ajWo2EdVCgUqo
TDv5qdkubWIGRreWxXlJs/sIzzWitJP6a924C0HWQKx6BEKLo2QBt23nH8C4wCL6yJa4LCWmpuMu
zR7JiQarIgI/E3QXUeQxO1MyVMiEdQqiu8VCp8DV3EjxCMtb39V/p82vN6tHjlVOLlOy7+JJgMN3
3+AiATPfv9ftu4tUFLbDJUW8nZLw/X5Vn2LRpzeS+2QVvQclHERx4oa//4ULOmUNpPjccRtsxd9B
h44wbbykbSVw03EVZ543UXysXHGq0RnU4dg6n6ARLIuFwEbMtsugHIhLYCXsfW8MPlvgY09iv0Vs
v+UKKEFVkSi3QKItCYa5rCO8BOWenps0LWADKzMBN5heO9+1MEjqlDPGNnqoa12UBQ7c4XNF/81N
C3TgWd5e+efPaJ0Ab/WdhHGMJPkrtlxrKIqf6UY/PUaqN2UJm7P/IRTblGN7HN+ODgyPRJMAdklk
IyJW+JKvNJZeKd8m+lv21KXadveDCQXMQfK2mdKo2I1tppOioVwuaUMPDNm8nRWTJZJmQtkT9Blp
Ijvx9xvfoQ6RCIILwSFAuSsQjzPeeYAmuGK0Rz5QtaSOnDU3ECzuxvQjgy5B1dI9QHktY8psz07d
9g/vsprnaWoL1APMOd69giD/RnVwJBPyqsXPMbtUGvtB5c8K5Mto8lhSrhbxfYlJhDVryrJfX7xn
LhyCO+waq45vMe0ImeS66edee2tRF2VLbmmjhVpe5/yQo6J5iqEdYM1iK0x6vJ0WBf3IGTzMi0mo
ObKL8mPufT7ZJaXRCKQxtJbfwAwMdLplUn5AU1ulj++kwCp9HCBmZqvNWTE73Iog9iSRRXJ1Gj+K
RSmcLAtFQwc9L/oC/Ca0Vc6ptBGufSOto4z2T/awxSLnZoEgI8PV6Vvv7pRsIJHgA431GNGRmo2i
in852un24E4wMcnhz//TaDKZ/PYSEMkwxJfUBEA1zmpOf0bQ7lGrY2QcvYgR5chyYUelY0HlvuKk
XP8d+tEKY+sX2qOCoP7J3BPOih2hkY0Esg1wuGFvQPxbLnAZAMP7gNWoShKI9NjQ79lwqYwI1T3/
uvCxxHdoQ3J3cGxIugGly3uQXCPiyhOPHHG1E3/AM8Fw0WcopNNu5aNgXhTMHlAcUCqI136i0dr2
t6imvri5qQ4XRoOv7YafoLpGSTL/hsgTy9fLKwFbg1cM2/GQFiRGPOVrz0tJEfvErSSYku6a0mYV
Zu9XyzeQI+y8XRC8C2bUAXFINq52YaOJ456pvTj890PIIv1Xpa0eNtQZ1Yjk3x3RTLwDm6OQc+fv
ev29wI2K/k83YaQPmYYxpURJC+55Xlul6g3cx7k2h6GttLgGo45rJW+579RKj9XjzrF533MF37nf
x7OrOqF/pz3jwalVt7iujeqSmxPgwlruCOt64YmwuKd6Ta/XpzpSiwVlaOZrTHV5KDrA/rKRCIr1
eLG1qJRC0ncPxFmY6Kz+h6b0BRjutsklnQ4OkEEiIrx9muoWRH6c7zm0aKmrCeR1yXRckF1m/t9V
T+fGAjPQdHQ5dzJEO/dp1++6ZiYA4x3ynTVOYORqmOp92zJJTvzrfy7j5C76eCjHuQYbOEFb54fj
JsUyPlDKdVg7tJ/kO73GVvMqH4MqbtqUwbjtBE0ImVRgUxvphiIXMeUHwh4SEgH2pXmmILLQ2ehS
qPZpgJPo5tgJ67LP2e9TT+dVfXof5tTBZ0iFOLm7WEf/W9JcPtoy9DBSVt/a4ijuLZ4xeE+r1EWx
RLA+qK85yp5Eg5o836z5IypUDnriQx4ud0iZ8B9nPlnVBxyfzww1Wbp2ZFhhLXuNRgsLKSzOvURd
lDNFm4CGKvMXlLpqYuiIkDq7EU0w1Fu4nXCNl+HJf1qof0uhy/lPUuNcQ38D5xilzabVF08C5bo5
aTTUwxTYPk487sZ+VYZNpZNk5+uMRhWIvU27yICWpCwzrjMVjg0BNtQgblnn4sSdhH9v7hdTq/vs
F0XLxPKpJ982GiQd7gKHOEIF7qe7PmlAkAS6j7Bpy0eo5P0pcXE7tN0P1I+ZWiIZCfODBMzFZOVF
bpaGsZHTdlICMR3KNUq6OEya8ybyne/rrfAcKvYvzoinhbDqPYZmg+oHWKUwcBscqbN0kKXg1eMS
A9iWlMXwqYSxopcswnOsQsp52hTbx5L6YH2DO8Nu8xN69xdf+P90r7zfWH4Y9qTWRlxCbOa0Ct6j
g5kiNmiRUtx9LN9wspzrB7sFEm3Bgy0CuXdo26NW7QPiNf1y35ZDihLOZWcaARpUQJbQ+cKDjmqv
1dY8jqA2mdwOQHoxsyJOQXEshPUpv8NQ9OHd7RzP1sIOxBoVmZqK/6ele4xo8OR759J6s3LoQ56q
PyUknRpRrMEmAdg9vT+NhiB0AMqMBcHfuFondCGNWZFA17GdtiEOi8DbSIo58RbUFed+arYRJq3c
jUY5cwJ9wUg6ozMSaudOz1sm7kWxCmjxsKKqox+YE/2ufLvL085uQYmRxOmvcxXnF9bigILw0I/q
xyt7OfZqJSRE3jmNyD9FjcgP0W6j9N+kU0V4EkiaguABporzUA5oT9AiGDgS0nk/Gakb4NjJKZeK
gEWKTNrNue9hq5xEfphfz/xEziwfqV7AlfdOuJXJTE2XfhynNdmowOlysatyUbdnVX+IEB8Id5vo
7Ur9mdHJBqe2bESTfft5XsbT1g1oj+XojwQN3nf/Pi8PkF2jRopcALBNW6AvcO4DmSayBnhOCXd4
su4SO9A+M4tO4jCtDotf3bmpR/iwLHuWHBYAIbAsXeCu2UInaR/8vZK9a+gXeGFBfXFM9n4CjxuL
Ku4+o/S/UF18lk+EuGbeHzpWcIyJzdmIXoQwJA/No9rch+0a5tT6ngT4/LUl4C2FKkAiMtxz1abS
VGEGcJvdwPHGPFe8uxqffmg5Zy5BpQmZ97x4IDOuVf/ZBG1p2MS5VkcimdFQ0H5t7Q0fecvpr+CZ
uSmu53jWABXY6qvVwVHD1efAfk+E5nWEH8yWtIxa6FFcXqZoHvnTxfLdPRtu3+8crv08YtqQUSxF
WnsUu91HHjgfuZEC180cKn1ptP6YcseBvpjLvXz0QM8W4OBNfT3mmCqvRiWpuHAUwAxlNPJokTiZ
dAC4OoD3idEWkRHc1xwCJjYf7IYE0bdOCqpl2oKPkT+WJew8J/Ec+U9S2l3y4MeWTIxx28JaFSWD
3mnDsVhobgqfYDObHMPN7A1TtdljHdSVe259LU2tFL/+URSkrYFFCScsPiOQ+RZbFUtDkBvTm88V
LGurgDRsI3QisIeuD5ZQxsZXulKtiSEkOJi8A663op+3eRCK2XgPvHZA5ZQR8oN/GN205C3SG62q
29i6bsyCA2zt42RcnAblQhAnIyaeto/kZq9W/3HinBW5fAszeD8TD34h3B1UDW2vwDjr7ZBvbl7y
QMkf0IEv7tL7ef8Fp/KrhLFmcqI6GNM4otlDnMYpRQ8FOBS7bcMpL3gGNa1+8qSPiwpPXeSOT7mQ
Q3gvgsxENJ2SJ4iXAfMEoGQKoLeVWQnJIUG/nehrddjmkdCDdz4l5B2UsfyjPArgeda1QcLYhI9D
Y3YHORtpQVR3rodN2tH1HSdt7qDkF0ODRt4LjBOjhTd5stolSwPBKkOzm4m13ZVHTa1RQ1edTzhz
fV82n1VTMf743f0mX//htycA99bnRGH20vhZ0lZlvVZP1yS0+b2V+9CDhV+PaNsoNHq4zkgfUEk0
EqgqTeNCZLZ1/juF+jQqM1SLHZEyDF7iuChXio47rPU/RuGbWnpwFvYOTNGZwkdhzNPu+L8tDD0t
5ghwVnONuRpA/LQ59F39x8g7nKSO2AG2JzbwfBWcDachj7fG7x7OGjMh9zBv+MF4HE5jtOyPPzka
ZYDSWh793Qt2nlQ8M9VUmXA9aezGgHrHkqXDc0Y2bn0UvOvlWCYV1w3eJR1qRwpnXwFuTn+6voq7
aS3x9YdgL3yTcpLjHtrkbvLfGinBudvOTWCN1xYDNTZmnMOk9lbCkQ1SuwoBP3vvU6TpDVj0M6ip
qhJ46WS8bUO1UwE2G0T8L6n8yapEBnEdBmadelmqdChYH3lp4aObWo9Mm018vL4Xtsu4pFuWupFn
JPATyRenQJRGIZbbfrCCMeVqvOla3qKXAUnqLY5hSfX7aQmdltgJOB5aYmf/PR7MQcZfW4TnmtFx
9Cjvj8Y2NWEVfDXjkcwTPm4AZjMqPTynApHmpAG9zUSdX/BG8Eb13a58d2ZBIZKpNl0PBaVt00Q8
EmPFAEhfNkGcG2HEzkhtbiXZsMMgx/cjgcuv7y/6JKzOzQsNvf6a2XRHyn02MbGhW4Mierk9oyBV
sM6iOLLNv+kM1hrHFOfynaXPsWXswmI1NHgczb0rdvpsyNQq+KuEl9IraJ/cPKeSXIIUgcn+Ik1U
M5qZimTNkWJ7o14wfTzdduzhVDZBURXLQUPyCJIobhqVmgjYUAGTZR2N2SWTk4bw7QDetrO+tvMu
cM9dDEPRO2tnwpben21+7Q5qoeZDhQJKUNKhI5GDuRoqv4EkVkcGKYdxxl2CF8lNocEaLSgIXaW7
aMbBZdPZYMbj9NLBTUfKz1UsSO+/uvcyW41fbi1nqtdKiqTG98zn+q/9+6l/ZBID5FmihJIAfDv7
knGRfbnT73eIl9agOjhFR12IwtOj0kq1+xArpCQlZNCHMclNqqvBFP42CopptFXStJYcJ93VPNCi
blBt4mG5R2iUilHMh3dlRGrjZh6s7oLTprSnqZh6Gu94RbyW9VvzoNhKZYjGndwqkGBCziQDAP7N
pTToQhWiJhRc5y1ltZPcBerKK0GodWojARQoEvq9Cn12sa5bdnih9NR1oUJzcBoEMVpsiXLam+XF
TYGURIjKtRbs/swUkt7fWWX6acA4ja1oVb6+bF4QT/p9krZa4s+6n0NYPUsC7GUlWUiNzlpJGLc7
nMuLKkn254QPEcV5iEhtV5CWCB7wJgAMkrhwvRwBOORT0LoIoKwuZjWyTgxnSxz379WaB2B1L0dT
177CqO0WmMci2rN3rHBRi+cZXdq8mcQVJ+ykzkTY1gYmOLvgjqSnJzwlvbzrOjFP8ryr0uHjeBlc
6bZGg3VNmai0niEJlahF/jcveM8qBvZ2h+6DG+rhGSyey/2Gi7a+Vn3auVopgPnT+32R89Na6hIU
0LQ4xN1rDFPWvVIJy2npRTRUFqN2DO7hl6fJlJqePzTeakRBzrWgVEb2P7iLt8wOJVMO8x0K2uHM
vt1y9lzThbpkVmNdXixO1N+yt/J64pXdmsymQAcuvBVjxmiAeiXodfaLbD12yw+E5QewgZLNMLsx
VBFFGvmly/UbI0vCzQnZ/M5CAGEb2ICDNic3RwnS6NcaEI2jh+Lb3AodMNtIW4OVnbzqW+eDPz7i
ofQLKsGLT2wc3gKHAO+Q/YdCKG0U6n3RCOZHLgKlOeTS1ofMwTwi01lDnc1taIKd5ILZB49d4ghC
h3KcxkcbABmngkCowi6iR7jqU/+QHzrDXtWVhyn3wMbPoyd/du51ZEkQkDUzZA7/vLyskJF13yG+
D5P86cgHMGqW70Ez/N5mwiD8tFZjJIj/Ccv1IqeLpDKysrnR0ssIL54R80xWkATdIcP1x2ccDeMP
tlSuivPStRFd0/RIT5mXavuafqJHuUwq6y+Vhxtz5Uvr1YkXW0U2T4TPTmj5r4d555o6irljgrPj
mjdxdIEF2ev8fX7Y8iJgWrZ7ldxAnIpvbQQ/CxJZ1MdURv67uB1z+MteAsJOUWFpLDPrnTFWJjNT
LbEBMVXJcCbsZzYyIcYnGT6hA8cIlW0/bXctOHOKVHL3nkeAXXTWzUzzhH5Y8ZGcBXs4ASU9/k2/
3cYRE/2l2nvM125bs0g/ukhEJhwKP4meAm/QjPhgRXJUJMewbH9oFUv9a9YSSwsVdbAPimV0yohF
c1CZ2oViRfjCooY7MLGMCtm+RrGgyN9XP/euXzmefOc4nL6rxRbITsAwLnoUT428THIiaaaGD3cf
tIOoNYSUfQYI4rLAF4wjt5SQgXKJJhyBOt3U2KDgUIVw02doOW/K4qOSQn6Cru3f4wa6jwi9plkj
0gpXPzfxwu6+fmuxJOOUBpdm6FO0BP+PLUJpV1QQYG30IoOOeeujhZoe0/SwN4Baf35BzjM8kucq
bWn6orIB1V55S2olGRWEuj82fHb5D2YfVayMCeVQmLFfr+UXADmnAlvuVyBX1EoeRBak2cQzLxxk
dC/xBPzL4LRfgFgjlG3lOEIhMyX4RNLSGlyAG43M6pyoYBEoYa3ajuKaXHrngYBa7aXv2WsQ3u+W
SCFluLwKcAuf7hzuosvNczIDHJ22YxaljiYf+mCdkViVlie6L5pWa7iy0RzVv01fmv91/GLxUQwO
ap0R2krANTG2TUPz5dWZDfz49k+YjO/e+01r+W9LiBSn16oOJGfNutQ+GIRyUdlhMSaFCoelvEiE
UaxvZrKJPPQXqaW9hBvNXMVwvJP6bKA7K7/B34a4/aMZLisjLjAFlvPPxQrPyBJeVV3BIzQm0/go
OdI/FetGHMeB3IF6yLiltroEE4YkAyKDdkc7hiMgTb9yKhDXfHg/pVpTyjXBxjA+kUJ2NwrSa+Bq
rb21xivzKYzCSsEz9c2nTQvuy3ZfQ1if7e0iI6lQmDhBKaLqyWOVsx/Wec8SqxgLUjW3ioOxggWv
4fOCPNrGqCnFnStlil/7WwqGGOp/bz4W+GCjIdtQnvD957+g3eRUhv+sFYxneqSotK3x96iQC5rK
k2KX8QcosvuPEo8hutM/oPkanzBTFWpFActxGdXlHNMU2vPmYgSFLZWnebPG/4oui9gXY9+lj6LJ
oA3mydW5fl+1U4n0hlKJoKxtkG9tXoIZW5ow20u3qYPWw+CaDuHb/DdtfvZP/hdrgFTh2HePot1C
NJcqTyRj22pK9mwG8707opFNkZJQL0n9RRCTNJvrFE5FY7QI2TaQVi4ArPdGFZ5p0SV79DST4Mcy
kxsZ9+AsTgvDhRQ9shct08o9c/lnIoNmPPYbmYivGwORzsN/UJH9vEvDu7FOMZ9kTzashLmy55KP
vOVn/3ZeKZ63qLQuUG/RtrlU6kYVF8h81dWotPZu0lkQYBbU24LmyTuvuYukYr/vizamzrdIZcb7
rhhxhkG0rpwMSnTVLKirMFZrN0X2JR5erRuZXsTAlroEX0F76xXwFfJBnmiCGsuR6KFydmG/cnOO
rlhDpjPVHdEnKmQrSzWAAs7mADWsXQKJN/2sbe6TXBOl2eI7uWSVx0eBRrbSRxSf1ghSeCxyQKtX
lAED0V6tCmNU9zNaCqn7wH3jLQeGdHIYX8y7Zdl53z5SJf0D5PSbZJ/31grW+3R6LlB+dx5KIriY
PJ+bxQ89N9hBl9I1oFhXwOxihWn+zR7ARUiARvWHRzSwrd0/dQHfLzWKQiSAf22amQY+EG8JJ5Vj
T/7UVdUEHmqRHEiP8VXs/6N9cf7/blanO+OYjPdsKySMUmDDH99gWZffJm0PC0d8FTP4dlygaOpQ
RXvRlKjLdy9kEw76lq5WqTRl3oMaxAcq9AxhR6eU4gWtbS3xrr1N5v9/7alcpmuKymZeLM6BIDqq
NdccLRJLnkz0pWJ3jjvzu8Yu9q6Txk+a+Y49hXhO+VNzkdwGsjbT3Yrox5idgpWUvbtP5q/yZrKT
oCaNpzgUHo+Gcp5/bRPpz9nRn2oZ+03K4vfVHk6IVUk5J9/fOisxUFAXM0aoRFsT77ru6kAQgKBI
o9ZhAbgeROrW7zE+3WkhvU3Ig/4RlkiiL1WsLtU6x4AajQr8ezVLHRwSyYrOL8B+Ypqyd5Ji91qF
O3M3oYObspmRkMuKcojSqzXGEu1QRX5Q0G3stSnYPUJ0Z5g23TPjeR2cTNH+QebV8Jr9bEuziB+9
mbj0ldqvFmlqNDQ+cLY3s+cl1o6keHfGxmIlefT1fvAZysNvj+00nmqKICLk9keDikX38tBBZ8Un
yRVwqklM5/akodXnFBc6M8XYsfwN+Clpbol31SGDJBQ9D3IVm/1bNfSre5bCwp2V9g0FSlmXLRnA
j0Z07166+p6BHjY+hJ7/e8WUa3RgXAa7xdIF0c/qHaYdqF0HJxFVBOLK7t4hCIEGSclJ/PxKiZZ7
orkAQkVPr6IRS4w/JGmhh2BPefCQbzxEXLeDWsf4CE4tQWFNFGZMtzLjq6dBC+G01/J2mAytRcsr
xKSbcrDTcjoHolbK5aimhUJLTbgJjVNzFCWBAWgnP/dxEKqgmYxWhUgUnFMQ2BNJzrBuzRqV36XG
VJ3T/0FRzillvsfmSoIAMH2PU+7cJv6VybQ71nYo3tEGXMKyHhrH/99a6wkF7Ypq5ZhMDjBQL2fu
2j4sKFeliTCMkCtnHhPfYztQIRJxAOf2wDeaBvmW/20DVOO1FlW+22xwbLJBbNp+l6Fq+XzNwOYa
cyGlTZ8GTFgBJEmi5gO7U96ZXZGajTSeRIx7BUI4QXW1XsYQd0JcZ8eNoO4gvzPjeeydON7w4N9U
DSFwsLMKg6bhm4bLKXg23LNfC7e+WhA2RDbtycBS3OV5JX2rhmhOsTVAR0/bxDFqBAGPevMwdapy
Ibp+03xpGNcb1Bg4tqPNlHzApWGWB+yB6biYqleMKERpsZfC4ZQVHtnUNbFR+iVoUOkI7W5txWBo
hxtHyRZlresW6vO4FJsNLIMECcV2QLvg8ZQPIvrzeNF63Zqny5brEPeHSGTzkV60qV3HdV2UiWtE
TxHHFz1+NFjNCEKyL0NJA7jKI9ZrUoCZZ4WxYSjb1YEMrRs5eN77c8X0kIaSPfC+Tqst0+Xo80E/
4ZGE5PetBahHxpFogckp74eT3K0ozHgl3VKrhKdy5USWZWnqWtaWtFqLxJoItLwI1FP0Ia/yGv//
pcgfbVs8Usg5gXk0AdPqAj2UOawsOtffcycWhT8vb1EjKji1643BBocFrONcr2yFgA1QmoA9150b
t8KPVg9pEJU9cOwlqGJUz4t9BDVafRS6Q8s7T+0QrG5atHToioeP+yFGovGueK7r6TwKClOlCaur
Mxum50QH0Wi2staMWruGcvDEa09PQf2YqJ/s0BYkcBrydYjvEPl6+XdmSn22jFETwqxKueWrroYR
LEiltWgvSndDCrkT4fBk167PLJsD9hmO8Bgi/XRGtZoWVpPnbfkhkXUPcto0alsjnYnImwXAFCjk
umBXTYqP3DmfJPzyTpRmD4ws7RMKM8UHlpFLRHkkIX64BsZE//JjHr7MmeoVy0GNRPlKkt3na1Xo
qumV2sD2jFVogIgaOdvEH9wmgrsapp8E8lW6rKDtYLqpNprd6XJT+7wSJVs9d32sDGE9JthyPvrW
6nXCaI93uaURI8Var27y96sFa/EjTP3FJ42HOBtF5A74b5sSMRLGYe2tIeugS8eY+xa/0XtZpqML
GhlYM+jP5uEwxV3J2N4xVrgcuwHxbBF+4CrHIwe8sYC2Qo6wwJmRWhsQPhIh2JOpQWLmO5+y88HH
cAPuH/wdsKAZU13oyhi67yupqc3/U9m2Yma0J/R+odavkpjgGWzfKJIfY+O26HqpFu2qBE6qr+u2
2M9cCJqrVU3kfzBwKimWhgLM16sqkvyRBOYfslUWsBsAseBx3RuvE/HEBJvfKkLsEgYNa6LMmE4L
g4E4W2XnFZOK8uEyY6AtKwoKd88v+kAdfjcN9JK5iHyo0QyWQNbmcsHX2W1okHdP8cMZ0Hl5udhm
srwXjVoeaalzTADUDBbdDI3R+1ew4dZR7Gfp90yqR2CbovywqiKTg1pB1fNacYbwKHUFEXYKziRh
oelk19iP13OTGsqPZnUmQ1iQYaWVPyrVm50skIB5ZFkMORxfYElOpFj7q8xfkazT5MoKXc8etWS+
QVk59O4M8szV+epZDQEYiqTtmNOssLQN7gAKWoDwh3PfFRJZL0X6wqqiroKK6liU63TB7VFSaya+
sxhHlWV5hjwdpS0n8K//z9wfeQ3UfV34rxA3st6eL+8ZayftZe4CxBq1dV+dGZDDC2cit0sqfPeG
iHUrKUO+c9LsFxqXR40SvGsAxksg/rVYkboy6/UhBdhqFCidX3Mr+nVzTzJYUkbdCTDg1JqW31ME
Pt6BnDeHtAa0zOmg/k3HChMASYUOxkZ+5LeXUcL/s6iLAL2JuiVRltGuePW16tYdOGir6tQzl8/t
yDXpoNmQPms7xrVPqpzWxnJf4imJgJU+nr9YeJeie66jdaouWUGIN9MZipP6okdp03J+qhyMnJuq
YCVqQuUJqJQ4xua7lXo1LlhVmMs2SSSFlTjkrIy/IUMOgoUvHsIzZUpSIyRaaKvjKPLqth4heZ1J
fF9SFPXf3pleavwZ1EcuP5UpYMybUmPRqmj4Vh8eUIHvlg09Y6Mg7Q1h8rEcrzVLQ+fi+ca8dyF5
dl8b/J1qMA8Fxd2JvuQtht+2PqCoti1DMvIdI/JLkmlGlo3ARL02uiv7iayRdsPBhsPoQkhVXcsK
FEPxKywDWIj003i69iwmk8hPlBTvgEmVdXuuBTna4zOtIe9uMAE9czELwbGDR4kKQ2gc+B2eY8jK
xKsyX+Nm13TRagByBLt+6ISCDpyXuP++L8mzwaWOsKcmSS7ifsrsstaFKSsRZ1CuudbdK+3jHr2I
NG8PsKkUowiW0ELNe0D2Oxn+o8v6L0ZgZifZgHkFYcCkrABytcrWHckrOgoLgD2svD5yF10+yb5V
1LyXYnfIR3OlPVJHdroIofUWNq6FPzKKffL/gaFoydVCLTrs6VYCco7yo+jGmUT4kf1UPHpprjQv
bjqlErwDPVlWG7czQHQUfEOYc9HG6SjET5Xen3opOjnDdJ31Tm1pZRQO+jikoiwKCX2LqX7Po5cw
XDPlyKsD1UcVypZ40i8EBmK8FjFw0qNnNf3GpHW54mM05WXLBSc96bmd6FnVcAtFi/cNdqIhJ2wK
jijwwoi86p3vAOMYWVmhP5reA1Fr21ev6OMc6TQ8sGgtcoFzOlIk4sH4Plz9lAavjLMY0cJzvCgO
b+SsWAXu0jX3b+uThoz5olidkqVbjZ07XIIODXMF03bO5XKuetZZM/dZaxInOE3QqagxkGtBN5CP
xi2H3oaR57doLp2H+FBsvBxN+X3/p8TQ47hxaWtC1/pUygCgY3rIupV7xnyL1Xpz/Xqq3Z67ZQAK
Iv4FpS3sTC21/pHvF7O1vF3t7ZiM5Gq7sv7Jhw9DtlzBJaTh5RLvyp7zBy6zPJEK2ACb46dfhNaA
K2PZ08Ui/AhTKm339R07bGCRHUx6IyiiNhDwwhRnEidYfVqdd3kYiZNQXIhvwYeh8o2FmQormI48
z1QjlcRsneX5HaHDd8FqMLWU3N4JBKPsoC62qFdFLX8MG0/oGW9syYc+ITtbJkfsc36F1gOui1zz
GzrMCwbsXn14+bJHiq9Z7zQrPdcc/NFcoLo0wLR5ojo8xaKmXRb4AE1MLURiJN5cib4A9Z+sbRSU
KjqAxwmTBTNnpZ52luPV6vbNC8o/JwsX9hIdGJsDVycws9CUl5jc0xQ8qgj2whPCIveEHjfkCjtj
4H4w5sLhzFJviDB8nsuOOzkCld2SGqkGK8BUPFpUdxHGU2vGQCMSD3PctsiBCNIxPmxXzWTGFo59
etiw12X6W0h008L1VSqrsQP2q3McZhyi9Lpq54gxbV3qKdWbAatlpgHKO1T6oQJdXep4Anq8Zc5N
6lp/N8AkH6kFbXqXhERQPspbcBmElAPMGnBPxoFskx8c/HW+9qGULwYyxN/9GW5J14wVwsQMyKpE
JAo/hacfpMqFnEZenTu5P9mmPN0ho5vdf+IZ/82URv9c97vO4fv4T5ZIjKT1T64dsVf/gY576pCb
XwPIkiY1cu3zFxE6WZ2akcuSCLF/YaaEYiocbPjqKwsRsSkykUk4KTWQNfg6X/EkFSgVl87u3q8C
t/OybdUztJAM4hmq46Rv22XJ+t4iGeHqW4XUWo3z3GQIAKsfAxZ5ASrT0m5Pre1mc9xB85JlNsVN
KhwNvrGdYQ0xT8pGGlc2pUrQJCk6RQsLao7wZJQMtaAindmHGf7uk6TbVTto0W5f5/6bPqhzc20+
Y3tihPp83TZAaEsaQFUg+X0idTNRZT0geYp6u7S2Z7wPkqOOK9PC2wntuhTuo+5pYpFTq01gHqHr
E2RiC154czoy21knCROVLBCcjWsPtE2hWcGXLlEF0lEplcInIQQglRJuNxZWCjmaIWVMIRMmzcyB
HksWK3t3+2cGIiWWrZYzWypnqkVC9Wu4uccFPa7zjYgT1GOZZTlTbaS3yHSRfuIj825Fv0ReIC9S
1+3Q00usX18Np0OJcrpJGzSHGwEbbWrz//RHLUwtkUF6TNWzRep1PuqwKnHEP/KsVC9e1Jy4av8t
8OUrH9vH0694J8eUeCpVzWixmy8SQLfPnczZMSBXvDYslnRjK86vbjoxp73zk3q7IYSVj8mu7KBW
hBXt3bmNbDx1firLQUlczfQNB5n+qCNdGexx8nLXpxZS94JJxg3BOzK1XgDRWd6cEbshR/vsDQS3
vHDNK7HI2BaKtvjjxC2HKYJLaTVS4+VJpsDS6pRfgZYQbDT8U+t9YkA6BDWnHtm2Te9pEDCEXstv
9Qabl44/02578qJCYlACfJ5oqyPqLxWYALqEPKlh6TVFhwkhWUMHgsyeBYmtzwstO2X523XFXWbw
R5Vp0HtgaaMfI3ghDq/pQvzTau6B/3GLEI6AZ2te1P3nMPeQdtRzyYyomRsobgsZRv4x7cpqzXri
P/lpHQrGUKQnrmR0V+dWk2nUuxf2HzFT+tJp5mmNhUZDwvX6gGndxqcy3EtSv5KL0SA35Tgmaeng
5T4iVGO+89sqQJH7X6BMRDzU9Vz+lCQf9xwmKzCvKb8PTNJCVlEWQW5khupEB2JX/4Jm8Cv6dNoP
89frdk6RCTxe8tsjD0f/myy50JutrgTzo8GNMPWFzr1734rKlzm4VVymiGSCd8DL4fopxEL8DM3G
iqcDNqSs/UsTt+9gmEvpx635Y8Cm7ziDAot0QnCYRSTxD8vOoTwwJZFzaCgGXJ6erec/4/EDwFPs
pKRzmGavJ9zX4JLftBjXMGkrPW9KQvi/XXIzEyoL9SeRINVeNOSzPEqO9PZ6ylZnNlBZJamGIC2c
1wONjNg6zSVeUYkrpVuVOhX1lKhwjIChH20EqKUVW6EBZ2fsNbaepNudaiczsleFW/QlcKlY6yAv
ytdcfJ+WGiIDgGBK0ma20wk63Yo4P3y9FgYU0eHjT/n5zZJt6UF3SECjQDLoYrnN9ZlkXjgaPhEc
TSnmQnIlVfUWLMzxaUARJA5soGXTFbhpmrZnbUzOtxw0YC7/HbuMOzxOc+r4SmM6lvWVxS5PL0UT
g8irIVdtkXTYx6ojqwxkzamLb21w6gDARciKn4GxUYkRrPzqj9FEoTk116m2ocrUVcP+GcMEyn+M
9VMWQB8tNUWKD7EfQB810zsG5rwR95+4L02QnL6fRp3B+e/kkswomseFSR9jV+9oaaRa7qvbys10
Ao86GxFqSEcB36iw8rFTOkVPFZjVa07+8LNhCDrKNaiSX+stUi2zTPU8qIxVs/Adh4DH2hND1C6g
/l4d80RFp6v84TSk4w0Qy56m/1AuMYiGV8D7YNMcMFZJGLEG7vz1eP6WQPZvKADKmE85AtRjeNMw
SW1YobOTW9mvp7UuhAshiDYAJoh/Lpggybw9OH+GM6PV4ySwj25Z02Z/JWzYzhFBDFwQb0HbIoBn
c1Zxed2FhVpusn3KGdMAUz/Ucyjp6aZ3iHl9r+p0U3ejbVZJwdaWWKmaqMp5xwSRN6Sbym9guKI5
cGis7aegpUddHMdm6VzgUh+sD6C/L7ugBcYHjL9tLkatQ+KL6dIDOxR6pUSnM+amoyfarYtIwrtd
jiep9JPW3gGVeCAJsnaohgDoSKrc/X26L7SmhfeQs/FY6Fw3jw5sMPGNWaM/hhLbLxct774IU/O2
U4QHRp9+hJhBzhjV+J4yOo0OISI3TuGAgVwpamuEt7o97j6nWkcWCtd6eMSWf/vQ04nNjZYhtNTC
+hhef/1rcWI1Eu7b0IIWVadNqykiBvnng/5lFGMEHeErb/0lSGwnh+2aHGQ1BK8tZsU4b54MJdM8
qHQ4Rb43aC/ZoIpoXnMIef4to9S7/v4bPi3+EX16vEb0FQ26mTHR6iERbAiNo0TZ5oi3GTb8dWx6
aePN2YMrw4pz6M6JiA7SaSrfyuCwy7R/o1B0LWb6wbPxBBf4Uo+oO1phDNm7fuM2FvA5OXZpiu1i
dlQ1V8g0GmYboSVmb3ICfWTAQAhkYIrd/1WgUganGJFs/SoV4bxC1g/E1KzVbjaks6XMWfxPrZtB
NR4UmnMfAha6Yf5VmC+GoKCK/gRV6zpT/PmE0cp2+5eAKpiEfMYYDboO6rwwE2b64Y/cR4SWbXkr
yAO0o64zKQNap9h1MvEuFlKpTplSQrE2aNGMGPhW0oSX8DwvtX8VdVeVJotVzKhyR+elDy1BG45r
jGis8/xDOy4q+3/F0FJBDMY7ZYGFqQi/i00aOPmG2Iw5mxchLsFAFKeGZFsLNveq+P43SyO45HCc
/fvOrMJi4b19896C7HV+fKmZTbnMyGN1117fYoB3qnqhG60miZN9b1TipNljAALKUdIDWDO3NThR
RdR+2QoF6JXlmbbYFrovh9CD0JkF5BuYTtCbrcAXtZvfwJkNYCfNUz9HDaDfKFv6iD5YBgxkuEmf
V5WpTdcQORVBM77cWRPYoCMwHng5WnFJi3OopEOp4wUkd9qG+JmPakwSV6RremyG4aaDrWIjKR0o
CboXK0IDcCGifPGB+ho3qLlq05zVMgTlQFT7YD1FEh41oIm1djnGCH//6al1G8YJc8OPYqth7+5S
bDwkY5xerZf/ZgAe8IpuH/jrCvls8c2YDLweLZC/OGOAdE/gwygo6xvtJvCTCRgwohz7LNhBcC9P
6PsyMSDhzN/wSwltVspA92c0x4Hzr0KyrK+NzmuxwBwwMOHtrN2YGI4Ncjupx2A/A/+JVMw5T4Iw
KR7wVVgOj21wSXFpgiUCMddUL22ef7LKshrmmSKpmTBnY/8mz5+v0RCxQLrH6x7ui6orOepQvK5H
SZFE7adli/uzCbbF5NY+djS3JZihopz4RhPoIRSCFCy0LVUS++r8nUmgXgAibeiLwBqUDpy9EXh8
FNlPReO0lbYRdtVHY2QLv2QMajLMZSmZ6hzJb2QCj5JYfdwEs0xOmn7HRcAD+ck6Mze8KuEsfaxi
1nqwsJfo+HYYzIxYh9dC1sB4aCE2Lo07mpNLEewEu7Je8FEkvfHZDTdjItufy/iWQwM7yLWDWh7t
+L0kpbw5P8X06wIvzTa5lavz2lahLEgFrF4VdLFkkzv5kSPKOwspg1RgPjhpLIGX9Ur1u42M2YWh
Jng0zwjLo1j75xRpC0289sekS6R1ZxHlJyPL4AEFN7vhPismwKOseqOBvKx0jXqm1s33VPcAuZN3
CGEjaAB1jG/KmovX4e47FuC76NCkvLwrrH566mLrQAjQFQoi+vKW8tGbpuiR+0KPNlDMd7tuXEYp
t5eOOvnFhAzvn2ESTon8OyKaxaZolVbn07EsIPEL1aZSgWR5UcX+k/QBv8TcxjNpn5Pz5UEZO77V
XVKO79xab+ervR0c73gnSFvASsGz++DWQwV8FAblt9ddqatOGy13B5//rSQ7VpvRZP/KTaiXGagr
wv5P91o9AcMMdEgSdOwJ9Wod5M62yKfUyxXcgu3rudVC8rb31hib29PiB4NS1y+sEsIObOBjT/h8
4fW1UrS2psOiEjCE0HlFLdRWsVE1OekGEuRto70LftHevYfR+vl+HZ+GSYY/0UWCvqFnyAh2PFLd
OtBQdjMEqUQpOQqYs+zdeXBnGhPMb2DkQMTBG/du740ZIQwQcQlwJAffGlriw5Ev2d2BW83z0bB0
EFG1vh4txnEP+K1NzEBOZkZsajHptPFQVlJ+Q35Ia2XIhW2XrD47HSEfW9JvEtOx7bDOtxPXE0kx
A77T0pbaudXHnvrbPtJhC0I5lNMDmMY6xa7lgMh1lfl+V8IhD3AEiFUjcL6t1PwdMZo7e7/cBJYF
dL7KZjzeYNtVVnep+j7trB0/1jxlhtzZC4MnNtXakre11QTDKdiWAcncm014sNNItcfzlCUNzi8M
JOn8CNYxLp5mlyboMz8CQv1SddJH23PWhIfli4T13C5GCzsCpLsPVaXhK/FXMRlhWM9a+5iXYpgj
zVPRGrsSsU5s6XRZcTmsi3G981Dhj9xLu8y5FL3pKWSaWwBmTnj6EiIUGKe+d2UDRpoj0PXGSM1X
3n/Potr3o5ApdpOyUW6tnT9yx4e60LGqrpXPCSCgZDCb6nbqqfiis7Puo5ANLPJnzRosfPzr/YHr
KVtfwGu3KMpHl8hBK7sotAmVtDytdd1/Yv9E2YgDiRlCVaKtktX7sqsrbhKAX9LGVetEdooGY+DK
yLy3Nc7vCTP5RKSV8J6NlMe4D6z9K3wULr/md0CSVAsNq1LaLYLmwbO4ZDoQ/ufFpdM98Wu/mjh3
alWOkDEBJBadBD54Lql8/n5nCAO67U7FEvs/+ytko3tFQf/Suarg0SNjptybMWo0H6hRmYl9SIYk
WvWTybZv0l33GWqhT1Jwn5IcllAuhkBy1mypd+YS3v+6Ab0I8DoY9nCKViJI4tqxVDgQxjkeSEGR
GYbenHTPpW3JkNaw7WytxUQk7Ie98z0IjjuevAaXOJXkyBx7lNntvYxjYjeR1+6vwxRdCk+2ins7
6hOjE6UYwU9j08Sq8f0faKeVFjTHxROq8WlO45Ol17pVXxEcdIpcVeUzFGd6//p3bnwiGTVl3wiv
ZoyX4pmDx26YDyYgQtseNQO1hA3sqEjbC6vt0AWRZxIZTyOQMlvyiUg11nJNzR0wWrgLjWI2mFAB
3oPXiBYzy3U8nnFmKxpMUE+9Ygs+SKhtIxgppCGWdmkQVt8ifCKl4JlirXq1Lllb54DaX/cL90ZM
K+e6ctxzRf6bMJbF8CT+0roQC03m58s95u/lczbq+Lp6/rFliilfI2SVjMHFvzY4TA5zq6uiDd+L
MwivpmEE9Gv8HtYI9WR/zhFcoVLJErvZY/E7YD4iS6R2FYSdd9TuhccGHrP3Vy/syYKM1/vV9mB0
Y3/lciSSjJyvQ/xnrH6cyylA24GpvAbNJBYhoiSOVdUsLEhW78iDQDTN5JSiNnv06+faz80LKXiJ
gOYy7HmvpxNzYyJxMIZLbwOT7YdyWWT1YWB7aLHTwD4y4AIdaXO1d4k1KWu0lNyroCJg3UGdSnQW
TEahBLdbX1FcSHjonruUAupZC3Bt2HanffC22LbmnpLTBYnrSS2Kt3NrXI8z9xZpBvtMmuQA9Rbq
dwgcOJM4I7dUH4aGMbrRNV+dBxAy7szaTgTZKwpPMzbkUpQ8Sgz09bYWQOkuaVG3SckJnSUfqCBH
dErQqVX9G23sH/+JvdZpce2MTmMdPPTV03SWt7X64gsatuquIfgtmaITgZVXdzqtl5wt5GciR9fz
W4OC3Xi158/egk6RjVStt5SemUJcbkMAk0Uak73ih4NKhDl/LaObaBLeup5Fo2JcUaeaN1OCTyTK
1ipabQCV9yutREdwOuxw5fLIpwvhwTxMonMDmnwbAQ4AcuMV0JxUjOvsYL79ARmmb+PctS7aLeZL
3EfEN52sdBuMxNHnVpwmPeEvKOJavl+8XGQ0JuwvKk6Srq2ZgdRDzClwQyRXD+4qg16pCs2lhH6+
FCdsFl99PYLCNrVXQM1PbL0QMkV3aNlyw+H83NE8ddP3Jt+c7SA5jm0pvPBtOZPbKOtRfVs9hz/r
dBiTSuz89d1iqlF/pSGQzH42x4MSxbMWECRZ4gD0mXWXKZuQh2kDgmVoKufDGITJ2FH0o0EjIDwJ
2cZzdkOGO6BMofb8NVYYp0DbWWFS8fs0tKSndVq0M5fHMdIaWotNZdMQxlqX+ExXQ024vcoXd8Er
NdFKnlE3PDVvbGO1JJ0MNtybr1zvtR8MPrNH5QEVOEKgcbNfj7ZxpPjAmP6UtI0DZsHNWeUvQ9yZ
Ih2oW5iefX3ScmVbWzyHCsrNijaDHY/c2DlNuhc8q86fqXimmXzpRGRmw1jnk+xzYf1wtVTETSEY
rPD+g9pwn0Ds0MCWdsfPdaz0lfFYItNgymThgUPEU6A42quhELV+w8oyaL03Upz2AqdowRCbdIFv
mSPoGdc4WMQqTKr/mujR24h8E7SNSlPnLRfCLZg+yf9sPZjc6tEZeH5ueNSECQ1X3hbHpBXva8JY
HVxhmRm0K0ziMWfdXYUSmT7OSddOFaUgXvK40PlhSl/uX7Ec/wjsTUXLTeUeMgIkSO51TxBaRveo
iixwz4BU/jOoibNodZtN4CrdESiMybMfAiJ7HP07XtGADFKBicg8YxxJq0VpVqoah2AYWnfRQ05A
9iksjqVHvnfVCVX/tT9C3ntgvuA3CmVCXm3chDCTAVe2mInPEv+EA0zEeKoev5hBpNTnRoQKjZ5o
ur78J26Q1rMCrflAbEdQ13BtDN0wgCLjzJXrMtw5SRMMdwfpKbhCvmApx+JQj5KklGYoGj1EfaxI
jsnJBSK/xp5OZOydCHJdmMGbveVudp+buy239x8LKWBgRaibginQZNLQIXQ30ghTpPR3nINUfh60
0Rx69bWy7B0/ZQjFsxyNUvJnO2T7IRvaaYSDSbIh4Dsg4bW4giTugyEqNbbxKZWzvm+Jiv55Z+YC
kZ/1vJ9xynLVe3ytRZ+0TUKZ1DutbcxM5qDi117LcYzGWHahvfDDduwDT1FUDtQkm95/xunURayp
c+An5DnR0KpKmpCwKiwTlMRObleRnWdq8pimo52GpY4fRFE5ulK26NBTQoIXoGEvRLVQBEZ0oXxt
w5Z/tJ3DfT02nURT4MxV2e+EMDL/GsoEJC2IL9KturYT621274L4IEN/xGndSXVnVhiVM6ow8L9Y
ype2C+LV4sonQUBqz4OCEUCXOg52VudJLC3ZxOkJZgmpAscf6CMt9knstJ1DXQUynV8OdWHUrRBt
WFPZdjBLGnuLkL5b+pGSGhNs3watG1gqZxY5Bb6tEa7UZzL5zpvKAJ2iDS31K8eeM617Jxs3WpqD
phu4zP5qNSJh4B+eNjO5WJ5gjHFWXtjOwIvYQGGlv0GZDwAAffEoUuPF0HQuWHR3hZp9fVTxUbgs
JPKL1RT6lXHT6ATpkNr2DTdhBNrUhVZvu3DFbDIYcSNN7jqDeoNqvRJNzU5voHXmXKrH9XKDZel+
YS6mXAAqZSCJcIoVeiLtXs6xtbeXiV9t4XJvNt+dY9OoWcisLE7Sv2vS4X79jdtumwHNbIV//Qfg
juusDAAODovtLItfLf5WYKLOCiwMq1zbUXHRSWt0i1N5j+PtDEdYG4qrITEQ8Mp9Y3Ze8/llwj8N
q02FtJ+o7RSF/7Pha1hE0qoPq/hTdeOcQxCj59w8/676vw2xYs3oKyOvy2AzB2ZEC+VugUrnFRTX
J6imvfQ7HkCk9YuyCf2yn5RA7NlK8YqPsB4AK/7t7HRAyv/XMsfgXu0hGHzzxUWxwz4CsvR/QPml
MeiAVld7wZb21OGrYgvhg9y6IoD3ZdnUtA5K58FERg82jr+p47/eqxkDrIpywUHhPVTcZPztaOkL
IdB4c7bidhd/Z5lU1UXgg6hp6FOK+eUZrTnElearE6XDIO1L12RsPqVOf5PCCilsDfZKdG/8z3VU
ViJYOxm1eFjhtqSqrYLglEpHke/37Q03HfIabkls5jZClY7+egiDYOrkL11fJ/szT//Hu5ayZ1zQ
NNwHbm3hL5pQd4J5ZXqkXDm5qLnTps/IdDOqyd51MAqksvNkeUU01eTF3FuYrqYgE5H5Zq/rwTrj
yQAz9BCf0q9y0qtrfS/L0qL48BxkGQ2l5zlJYHwiLUlCLvZTrNpPh98oSDI3JegFyYFdExYgdeCZ
BfpUso2XqC7xAh3Jp7W6+kRqhbf5CfL3QLkrvQ+FS4Kb+r7GaroG3ALdDUuvYNyoHZgPNdCqc7yQ
7kOWC6z7zIDEzEojLwjXDIRvClk9SF51yL/7N3fCchtwzFpCJ2egXm5n5vM9EXDwG3ksD/megHyP
nobmO4HckS7d3not8rqsx6ue0D8wrkCpV19lD/iZFYQuJbYRDgdGn8+vs4Ztz2Vvp9Q9nEdwqct7
9U41bKiT/cRyvVO152bQL5cJs6lETk0D1caw6sAAC2w0Eun1vCYSgvWwzlk0XWEtS4v6RtLQxbTF
CUVMkakYmVkQ9IW+5vQzTvg81c/OaieneA1bjKvE0YkLDlncgaSyaOzV0Mh/at4m+njNf1k+H3sS
6nWcxSWioQ8jS0/0w2D5XCoIqv0/SbGbOvw8qGf8SaJtbnSxmzwtb8qkYrU7TTeg/rjMkKlvcmxG
07RKqCxd1iIT5pgxrmZIOuSQewZ5NOakKzU5S2TkYFZibzQogzykTCA/l5W0c+dFyyG/BBFLzEMB
2jxhZF7ZfH2G7Xduxm5RpACfKKiVfRusTMMMvwufLR4wX1yQG2tNv4rOnzZqqPbJxB+m6TOpXc99
IKAOwFS8PaBCJcMf8B+HZGwBiipw5+qvYZ6ssN0kjp/vuNM4QR/rGrQNe+jKw0eXij4YNQVythZX
QNdAc6vQ2Ml9grzCRVmKdUDeBpy9P0s57Cs/owf71TQFI/0No4iF8ptXS7b3IDKlcXFCZk7kJoQu
oyfi6wA5b4eCnK7AAkF5OiH+Ka6XfBKs2CPdM5ZpVnetQzgYjId790Xh8E3Cd82mfYQ+A2a3ZwCP
Hxakiodh6zByBD2eqSEy2He/n+M3JSwM1WrXmJHmZxfiHe3ga8hReuKtZ1/0Ue9gGtaXtI0D0E3i
gZpiE9K9AlMpuOaKpph/p6dbFcaCk+2BGHK46JN+ODAmv/YbuFEpzfDDpSX1Yh4GeAmKkHi4E1b0
uKuaH0gnuuZubDvBrx2O6YwiTvQBIke1L0Jaa0EfMAU2lle+yn+SJW7Ry4FoFEmSzpuokAYmKPd4
wFhzJ8WwKxpzs1gATqxWh+8Q3+KqremfCHNMczjh+X2LLQ3jQendhlkMzSYh9fJgOBaL2Ifi1Gfl
LZlol9Im+qsjlJut/2nUcCs3m4MlBN7QFXQgmLMLt1BDti+uiAwY/oi194WVkqKgSoaqhQyliyrP
tBZWxaV8vy1ef+d7GTWlU7r6LhOpNQPgB6oawxudm82si2K9LOb7xAw8qMZz/HgMdDgixyw+TyyL
HpOOIlOjzce1bMsk/KzIGnnDC0ajgr0GAj3G3CDk330JlP9kju3LGBhM8Ce90H+IbzdNCFfaVt1G
EjOo/gS44iE9SOMG6TCFZuA5LTT8i4crM+GbcuAIst6/11GNcEbWVgqZzXqNPG5GZBAGcWBmS4+Y
5Tuh+ovj0z5WyzHe94FoeNZbLKOUO81ECEce++mqwgZso6/YyL76qw/p1ZP+P8+qpMBP54f+rH/6
oSJ20+szCC7zpd270Anhear2XPqhBVg3HWH6J7+rr6hMYc5yzeYfdfILoQ3S++3raxP+Geh6aRW0
uDaDlq6FtlkInPNJ9XHlxcSF3RPItp5jCQWAHFxQRSFinXgrTfBn+1QPuf9um8YlpOlTtrBbqrQ0
3Jich2lNL3amt2lxy/T96u/1KJjQyXQCIjnvB8FMiY1TPTAlfI+FOQ7tLRlPh5FMhWL/tacISraV
BAWiRsYwV0Dlzjs3zFHhZSyNpSyzkkYwhDTaTxbaCGSrLuVwOi3khql9PSsckWpg54guMngfl6QM
klSws2aMG0C9m4KIeCfiPt2AFV8265lzbviPbiFrfyBrxe1yTd83uJjTcz3RimGkYKocTvpWoRIt
uWiVaedQxCAz2kPLG/7L+Dxfsand0QLCPLa2kIUalVfnnjqVqlrljq2MO7B3PDypGMGXSa4bdBpB
nV9hXod9YVcXcintoYr/TE+KPYTShn0fOfW+RESt7r3bvRdy6VrF6bOfPAIZsDtIKm4Ynlhc0xpS
KmObclw87/vGpYeABAWK8CBSfkXdAs6bafK8o0+rFW6q2xa8O+nLKnZ2mK0DBaJh8D78G+0V0cnx
v5Ady6NQTjFa+HZzRF+eE20rd2fGgsWI/wFvu+/3Lgy0/5V6AjPytiLmRAhKWTvOjeQNkGpbweMT
hSOFD4jbFcGlW4c+cHU1TU9HYmu7KFi7Jw5pHGHeKulZkq/etBtTut2HXZcQpFPhfOrsnOjdGQzw
8KjFtgVn0azyzMZ6PW7BUF1CGd/BrJUUU/lf30SF2txgoxe+W+JIBigqacIvQ7EhXW8+dNoSRf/U
rkbDi5CqexxLERqBjJCuS/CHAkpoIKpUFUUUwLgGb0LMBsqCf8aHkfsVxKkUD0sbii3hHAvx4W8s
eidwcAB+8jfa0NiqUmiuJdPC1WT+JP/ontDxCYamOuQGmtpBnbwL5SrGIh2z7eaq3n46obS5Il3h
5Sgvqd4Kk4+CrzWr3BGouN3S/bWgZSVilPweSpsaUMyhTgGVcadlamtlc8xbMyjgDcKuxUZ3jgRZ
nxBRpMS5NcSe1zgcmIdKvCT6heKuOiG7mAio2yrXwDCRYMfTPF3+NkY8Hb9o3QpUPeBkpnCBHiIs
bS1YhZfRUlpXMto3YcqaAkySmx52Xky03yA5CzQy18s+AzdRHz2s0jIOLoWjM0zMc6qB9rZXFUux
w35u9wyGiyx89CZPoeo41R2ax5sbiSBv7a1RMhDV3nBEpb6NisQJd8Zq+hqWTOKuTsmilrAWE38Z
cV7aVzbuMcouau+dESV6duF73HIP1+pA0P570jfUlOKHYWF+Ba44vUhSutNhhL089dStwz7CXz13
K74QKfFNtcln/sJqNSLguJelmC7P9s3N+7vEGFJmnXEAvDOR9kyzoBKmOxF+HDNsDOOuwK03tFEt
yM7r/z9fmV5NcxlFjMgH3Zm+L4cJqds0QmWGVksewHezCgdZWAv5EoEoI2fRqxv343BZSlIvUuiL
Y2M7qX7LeitXUZYuBdnGLAjMRTjgONT8dTO9GmgEks/rkgJeBbwo8u9saar/8TYqEzHN2zuPygxR
7pEgQxYx/FUWcmsqSlrokhGZM+a1SQCs60u2WgacYews1QvV8B3YS8F3W6UlzsSkWyifE11bIn9A
1BZB6roMvuqhz2EKYi7D+gRZE1I4Ud0LCmtDYa8eH4LyJuar5dXlisk7BSrde4Jb9bzQfI0D9+Dz
FQzorh/D4GfIYuJTVClfeTTA0Jc4lFk8TSOVnSW/NJA+fkrnY33sbAYs9bu0JhvV1sRZkFC09Pmm
AnCxA61kETevVFiU8oTQgDGtzIqzeHn0rkV8pFZ38OBSaqcNyaK5HLPtHmiVHSzBRxbDzAL9Ljpf
i/nk4WnyD625QiXDuMe77mfrbyOyQ53UdgErY7XqUjWrAPmDCbX7qoy8LFI1vcJsg9E4mukZ8+Yp
YrLBXS4pDH7CT9NuPEi2fYjIsdjE5rtkMKvpPwPSgaYRW6GSkwfG0xmHuUrwGfrnX3uVbco0pW/m
sUAQrZBVtOYMlxpQtnf8BamDVPvCMwZrCD17vcV5HSw/9u6ZPAlZL8hR1SC+v4An3WO/Vi7BvYxv
825EQZlpBPKffbTYx1JF+UIl9MkBgJcd9ArxKMsuGF5Ztq2QVY1ibv5RcO84V+dLHMtMJ1j60Bms
nQPRVUKloAksS1CnUaVRFePyLFS8xqyyYNdqavNw4iYqJOrKfaw4f+ZtGsEcMmuQ1GDsPmP30BfH
pHQ/TDEZU3N0hmlpd+33KFgTWzVCoLTj2SBlZA44cLK3JtHYkPGF/siOH/y9S796I7k1VO4zdv/Y
NLTxJNwZSujJHcF+CvfzCvp1f49tXjRFNIH2qEA9oMbyaBFwjyE+uRW7fAe91GPba3M8nWqKCgoH
+8xksCDLGxol+veBZm6gScrM0+llEinwN+dJ31jklhlRffMrC4HWUq4SQ1Y1lotEhlYgKvtVNDhY
AqPCPPiy0ktrqcPQtRZswve1DpbQx0h+Bll2oXisd8+cDgXmA6nFrAoW/ElsIN8+VGlt3wTUkn+c
6Q+3YCw1qqZBdLjv8A77yhymSEXRADmG+GzfFeU8u+2FLESI5o0fhdeEAInZRlI7ZLDVJxcBWsNF
/fQVOt/o++zxm+g+ZT5AmeIFq5guQkRDlT4YapIGj7TohrHUZvkjGUaIiLWf2V5IcDoy30yuLUwQ
1vhzxfwPtlLKc410mjvC1NU+U5FxJudm3H8M8+8iE1Ag4zrfA8xyy03AUa8O9EKu99CILAmugR8f
b3tPmMstoyIQ3GlV/1l/e8mqkbDmctq9gyXKD1FlaEs09bTozosU90jFBb0m4CpW0CzX4dstjXGk
BdiohN0qEYhEE/aZR80PUmJYuQxFzcgKwuIgWg5cHCZNtaw9CFhme/ct87q1iqYair8734znnMmT
sCOpRPgwG9cLP/u1ketCOxJwQNgk0aWL6MvrReS14PHGRo2uVC6D4duZcXnh7cQMyuAlBZ+kq1W1
xAgLXUwX6/g0Krz3XY0NC+nl/x0rI+3wLh+ZzXzOzxYpcgeUUMRuIukZTezB6n75pXSXBQ/9/4MU
FbdUgVmttt//0vCiFeG/BbbjpwPav8/+dLjzO1BE/AKiDf1vx9zkz4pYx6+ijY/3Vd3f5oSQCiJK
SK1bhLXfCbBKVRcAD5AjEaPgqdcIjFS1K6p2SylurtwhyCvSZCoBbPN81zj4vWixWvczhWVY6Ebd
GynMw3D9iHCPgS1fzgOQcxoH867cWBstBkevsBDV3TSoF/D0xSQUWxheZr4XNzzGgiSg2o/8dK7C
v2Ui1RViIoseZCAzWPGskvFBxta6XSvH7SeLBMXZfGUc7KoHf8zQQz4d1h1OgYq4nMKYuCLi+K4J
EpxoJFBnROaVfax9LgEc1cS11HShlaoPrtKYw8iVcnvjiamH0Y70HR6lhkJq5f4QbDLkj5A2XmNt
0EORgMF06O+7TMkhPHbrKBnAukSNbfv2jsvngvD4P12BSEVq9Lq/D2X6S7ap1UNN1NsUqUYgCgJn
BTx+Xj7q3D7LVp36WsVYL/hxj2ZqWiJRftCOAGgv/DD+oaeKoG+hT20ZwCkD4VaHT4nLkujmok95
cmIUa2+OtKxOzrquoz+Sm9SzCFivK8RWeIKCqVtNbO9zydL4U/I3/tYokKkEMzp91o+XzAiwq4/D
E2o81qpLEoq56GG5SZ4BfWdT9mTsMqeHx8UVPajfCl8oRscF/6YgHJhMW+94aQiPUMYgSTsbKm7X
O7P5CYylGf0i+Oh5ozrhB8z1A3fM0JNzELLnfll+QxdA3zO28264RcE5115+9oTDSYco4FlJEzwW
DczL54r1zfn5gtA/xtAOxU9AqfeTSxRf6wP/+89VRQfTWFKlRCVRbQfGFIu9qI/uqGzoP5DPzvji
JTtyTpuRQAOJCNhR58rusm0K9oRU13Gp6GT3oFn/0TKl45jxq8S8f1vSCy6bwZe8B11s7MXXJf1Y
Y2QGrUnjjWpwgXmfkqTKj/gTaCktER4Bxi2h91J1O3seAlA3pszj1Ac6Jn/R2MmsB12yUVNbw5MS
tWRnzEekivOoSuGp0EaIWOnGOJ+pLT3+1sC9mJwcpxtAbPgbTYgsmwBzK4Ot9gqy2rIJJBxfbjoB
yuKx2HLa2lkZqll+xOZDc1bQN5DJvA4VlKXF/YoD6K6F4PMxoZwvovORRlJKK+GEfy2EyC9MUP2q
YDNYG9ugZsiXKq8JE3iy+Kf5XsNX5Ozezy/dpQe0TFzlDoVZUodf1d8JxnXH4FvaaG8rBZL0Ex0G
vrJ4n3mHe/+jpvgRkodthePuKBl6O6d8HPuKUiSzOMSPclRLTVIdvA2518uOGdp1YRbhDfMb9GR4
/f4n2GfmK+2TlZhN8fa+itCW/hgaFQHIItcyMwbhpx24acklCEWpFdnTS4dh6syPOAhsD3cYjcdn
EL+nvWdSHvlPNiMzHvboAtXKJZYLVNsHJxf+IcSjeT+Hq/mU3lwyrobjXpoxTfwxX33KND7EJQnh
rs3TKQ2mjn87Fxm4BVH+ms+cav9Iq/71Wc7BqJdd/WDB0IJcaxW8seU4U9y9Ui/oK9aTPpApbiV8
iQcZh71OCG8i/ItJoOQe2LBawxI7q/LDAOy1TtfoMC+fHHnoJdGywT6zAFq6I+lUS1uDhSgu5ON3
HD3LVWn8Iom/OYqQN2YnbUM3Bbqr+Pni3WYzoYuHEI/8iWGVlUNlNeMZazV9D6T76K8kGxZyBaL4
XuRwXbiffPFdQntT78Rd9uro++drHypyUjXh+i035pgz7LXB5aNGpY/9msBYe5z7EFXTuun9DOCN
bFPHu64wpHqYO7d6W7PABX/6zZIFq93OlVVnOOU6aAqPWrIYFDvWCt/6pITJ3BO6b+/+108LwxaS
z7EBMh8RAjywWtxU5hqkVEpyq3AMwUdiHoWAVfnJwzutLZ7ikKzm+WsSOsfv6oethLA4ltonO4nc
tK6u+6A+itSXZiU+09DKjvOFwKqnr843byPr4fKsUW8srq4Awz7ysYRCyGP7M5emKnXAMCaAvpnD
ztfqYN2zydZOFdr7mnHxR7F0OqOEpI36oGqY/wvFzaZv6CPn1ILgZPavL644OFsmebsqsImzPG0J
EXwbSO1JNp6m+itVnHNfRpVXuWM9f8uzO9sPLVDHAcflmS4iFAeW5phQ0nNec5uDeFRJPWdvmJKE
ItV2s6Es7DMLpfLavC18q7BDVLEl6DNn8A+vW1phb4DepelwkkBVCpu7mLhwA91iXYF9uUVdugFO
v2PENdlJHqPJMRMwYgi5vlm39bj9Z6ACCOpPB91OmSo9ukZPrmuSujULcJtEhLm1dFN/eEVOyGyX
QsfQKukqB85K8DdoyWHar5nAIYHvD/y64HlOAiJIvbfiMqukGpQBhI2i8pMaGCZJQGwIrOmDQKsk
tnWvpVLipO1zRNGYzCKx0OOU2jB6s+xOleMUZ8F5zMBq/TrlHsALa68ZlxCkLubtlMIuzJyc6omk
SUxehFFOd1HfWfraunORPuTeO8wzC7Y25JfhXwl+sOPn6dECmLfj22j2tXeSk2sXqg77T6treJ7x
otTow/ZlVDvcXjWAhRDkt+v6GloKpaRAGgQo5kBb+JiQJdsDITPzaBbBCTzebQQPsx1MdTU8t2ym
HCLGu48RfH/tavMhtHPowjxM+3BZ6bNdrWiaoIlWsZbONzwHIAIx/sn7h1Ybh3c7NgEk233wmnUG
IF8KsZTdeKWX6tT4XaA5hWZ5EnrnAdekEJJehVxWTrhPNQhqPAWTdkORZ4BlZ4PEGUppejnDhoSA
uuiAsS4oYC5hvjaKlf/PvlgOvlUpvaWNoS9mdqzXMNaFYNMsS3vzXmd4VOot1R0UXbJkHbks2+ay
OY/GI9QWCTjsyyunN4B/2B+GkceCf4OC0TxsO6oBv9hvRznadHYdmnKKGwaLD+6aAez6kH+bw+fy
41JEkiYrRh4bEl69BtEpk9Z6gsMoumBy5Mm7Mup6/bc2VQJH71RuzXtIWB7XKOdCc56fQWHPoIG/
mco57T4+faPW0zjpyjnZov0sZljIMSsaS+5+HIoh8bK9iye6wI0hSGo6kYNdmZgjiluZvFW8O+yB
tIoXbgFwsIgwH5VDHMgFkGoVWRYU32SMZ7EUH8FDPL93Cto3DHSLghadHOioUUy02TqeqQLRhSBH
Kj2n4Hcex4Mjh/2gXt4r/Q6JbfqXZHJIcLZIp7eq6GmraAimt1VKQ2t1yt7DwyzvNX1kS2YOELIK
E1aR4HClCE8QcuADvLacyXjo9eplniidasTSkVJDGvhClfwR44EzmQXTCBuXSlWHW00qGJSIdYTa
VARabS1DJrrZ/1zyyhk32qClep28jv/6IOxO6QKNBSSw8qEbXj+JslaQO5iKcS7XmuQt27Jnk+rC
clnmAlKZVs5ZikBJ0LVYvgrftikMUKJyHwWDBs8O6xwqFENsHIk86YNTyi12iCWxSFY4feKwlm85
0bvYldJudE5O4XWIk0P/i1bJ95aup0Awk9UkGLqgnz1l1rFhtM7CCw2c1BEqRjQGhhKloQfegAGY
mYsn4G2u+TJYWSrW64BzrR46Um4zJN9Y1y8klp9lJWJoxDuG9LXabWvXTcKYOyqFaXQsyFD5ds38
7zcEXKhulPbtvSD3RBSwrbXiAT2yh0Z4TNUb0hmXjdx1sRbqfFVoiO3ifqrrFxnZY4h8c1NpGj4m
APe6g2LBFOV3KwyTOK35VKilrEW7+A+TGWsFCtoyIQAXAkHs6D9pkS1hLMvy2B+WWgO744lFQzUP
wVDB19LphcyRdjBRzqoJ9f/5styNH3dYt/zVOaUxhzZgwvSENdNwWilP8kmPp9CyqX+TqBFPg0wP
nK+XOzLy78BUt4NOsO3MKctwDPzqAyUXzVK4rVs8iwX/ggPVKuk759JTxvlk2xy0j0/R10UoceLq
KmuK5/dSBhG9u/L969vNpqjn2+OG5kPfYCrwgYRGbMuICPbHQ4lDDDKZoKKvYQd7qoerJtAdkn6s
0dz8i5F1gUzYnPagsVJQ2dIlMlrtyAnZEgU/kbDiD28H1JM0x+yRBqRa45apUCTh4Umeicuav4ab
PXF5mqxQknaQOko7vPwhHR4F6jG3w25dScoPryUunQaeap3RktT2vbSwWBho8WIPEAneb9UDldZP
M1pHZLLs63WlGdpH3dDJufnaKiHPUaY9YOi/gN8yUoPmcKcXX0pZtuSt/yuwEG+8787fveq+toBv
kJiQGPjG/9C9tGj0vcOqldP8d8mK/2nNCfV6dhSsqrPHQ9cwmwUk1mdn9a1oN8zi2y5g5Zd2GUPH
7rHMGzmuENc7bIkiWDfH0GkkgyWD4HkEQA5JbaEtXdsdMPDBPPOaRS+6GNStkn0wXAC27/pk8vLd
1eM0Cbs9affMbA15FxEL2jiLDJqjcC0ni0MiS8UKl17kHN/eQp1CZkxJrBtZVEa4hgNUq/gDll2T
VoFhRHj7qrVj0FghLnClH/TFAwNvW7AN3KDwr1dhTdDTBl0aq1Cx3p37/1FCK15hFTXJ9WDiL64T
OGnC3iAZvVsBLQ86LWbhJe1nNOnJmLLSIt12sOLYv/lIEFlLLduTeOYaYwHH4/A3tbw1u8cthkOE
EnXgmW+WRVntYxL3OtjpK01qCR38/u2kOQypThYE3Ria8pfd/daeld+sY59f3W/OAFf31d3feMt0
2K6Fn5PG/6KAcV5lw/LSadx1dSHTBpJN8jIi/UrpOHqEFc+TaIFSNSTzbr+CMAMIx8/o5vM9NDMv
LYJY3d+5X3Quf6tjWwQKUzKadxH7QzHP6nVC1kaMkJAfVK1Z8YpSMqSiO3Hhr2tm9Q5wBuBPxm4K
gZi3d6NyXm6JBM315l+XQhncyMX9m2zHVjNrL1K+ccBjfoKtjj4T2VWDy66Zrzan0FPQJKreSLxK
Xy8yEhIUUS+4LmQd+Qi0FKp9OpgkVSWNzsO3Pe03rzUWUStf0HB/2e6LQL1vjuqey4oP4UuWiC2E
7Y1PZ2pgaIU/W9pXiHqV5LBYsWmG8qL3hOMjMwjkZIeeOhTtZiq5MLOctRFPzCt5Y5aAO5h6tAYf
WK3FKnE4ooOfpPlXqp5xD3nIYnVMnapWOGMvbFIsfyUQ2tnFlWfZ2eCvVq2jylCpJ/iYrGbccerW
/yzvaX7xDsdNmN9XrMN6ETVGIQxTpsXAdi+95LwU6xFbJnvNjEYqMSBoUlEut5ptugUdT1SaTc4f
0/AENxbjv3nL1W0F+eNG+AyF66f+gXnYwsi5ibm7gux8S5r/y23cbq04Gz3ruc7QbTm9iYRUj9da
HH3V6I+zqXdDN5OjE8u17CdQ936s9NCup9K2cLEFB5TcI8GztscfYUg31Rbnedt1f5OEqh8jnQ5e
cfR8dmK4QQekotIcgdPC/lU+UTQxKxVXUfeDCp7q3/PdkCJc/KM4oMeyjglFKF1Gexnt6tW/VCY9
CWdlVqFk9BU6rtL6B7vIOqQJYZBeWyzUKYAd9KsNoVH6+tEpv4uEVjtw5T1bbyMDmNmNWk0mllDM
yhCSYm2KfnzukOOoJyncRihWx8wf0Us3jukmVSDXbiQSbe+Fc2RVlZFh+C090SvSvXd6gHQcghYc
naBEZW9kaXzRgEEbxr02ysT2KBl1AZnEpyscwBSw1vryv9JMuzb8t6LIMwVE4yU8KW7WWTVUDezv
qhbUPL+9cG7+/i4msThMpVw8xBXqUrLG0bXGh8tIp0kEcEtwvEYZIMDxbCLMv4nVIK/yK8WWXadO
DcVoNholLp6wZ7S9y/71lhZUgj3Cq9Bfj/5V672Z3nPsAF+KwTMDqL4aMz4JDtUacaiO1GMfR/DJ
GTXLIR5tecXSJ6F+my51qB2lwWCyx9PLF3rpx1R0EndxvDre63qJpKutFazXvuJ/FVJWk/czCalA
xaOCr+2UnUm8LxpO+dzu6ty6UryOcLnb6P3N0rX6TmoonN9YR0j/YelDKQbEIWYFnqEoQG6Hd5wh
Gb0L0C2hgtJsbovU82QnyFLMLXXiqK6G9q86QfShtFl3JVA7LBQj30nugdD1bckdlYo9+KVXAfzz
qqkQoTqBCIEPmLVt7wfIki1ChpGpjX9RIOP8m/oOxC4Vc/CBD7FcTC+IgtH3cwXG3ITsIbt+LPQy
b9pQBQ4vmiVCPuhfa/L+Jk3EtW41DYRX7j74HmbC72vNdUrpzqU9SnDDeq3efoT3aX/zLBdkr2/d
iqpcOX1fxbGcaxPynvbHMrpkZ2FVCDeY43pA+rAp4hMY7ILnGzYaYfED1BP87bDwE7W/fC2eH7fe
+tIE60ghq66r0hsNR3li9QpqhP0zrcHChVkDll1dM/J+US0olSJgiuPJYspAKBcedrE3PMCo4u94
HjY67CyWhXs9M1jpO07L5po1SAPJqK7CRpezvjNrFoo46r9YIYO4M/qgUsw2P+0HFUieufaqi+bf
II8whiF5CqHlcsztlhvo+0ldz0pqNOjqXpYwMhjzu5ELDk3pTjrpuuIsR1lN9CzeHBfLu47ykmBL
ZH8j5e9LiO9kap7KkKp9Bwh5Qiqs4d/5vaYGp4TdXG5MuAp1GujmR2wPzezMs+9Pq0mEQgsVXTUV
goMN8tQGZY1EFqqvpPR+fKBn5+uHkuA5lyY3o8pDiE6hhW1iXaQytk1l+PFxLPQI6GhtDVapLbLy
S2m3ONfpUYyEIReDOT+TL/+AWWThVjUiOxrrMEeY0370hfkF5BNIhre4kHj6aCzhGRcjAqgz2bkl
1W9jsUJi860uyZUh0MxMpNhJh5wxQLZ3tXuWXsIvaNlv2Aq1Vbc3gbBAi8nrRT29OnkxAQIINI6d
J/OcO2VOzi2vtKKdnfmxJPAHqn+YbdUd1UepUESJrZcDln5ZkpL+FXNtqSgBWNhKFJVRPGj6VEq9
2a5alhKzZAByu1goUu4Wd5ArqIwnnP6X2TC75OJh/aEfXVXhrmxluTIUc+uBskSr3TEnrYwu9BBX
exNPuzJHJibkgw98xKKi+KBkhQ0lrHzdZRlxxs/T3ojWDO4P/UOIS70b58wcqfvkz7Si59tcmAPm
Qo5skb1+mhdLI32lZ9BYFXPuKEwY8fOumCzsrs2lvCCRohGUuzaPil/3F/vSlMXtISUg9NIczmiE
UECn8x0Mn2rwSkfW5am8+ykReASsHOLn5hfoVCW6960QLpDPpQ5O7DiVUKkknBEUT8UCggqPknIx
yWoxq70c33pIw6ENPjxdcrR25IqYtZaGJvmjAkDyU/KLTPwBkxFnTT19cum+ZOFIEfpA7IRhCvGR
eWo00tMYQqOxw62c5jz5VgkZqBTeQCrejjQ9VQNeP/89IzsEL/MgJPxID/V9JFM/rrHEpwWBbyz1
60UE1ZbxxFg9620nu+HGpVX2XcRoH1l9q6wrEBDoVOEHauWMS9u8+gyg7R3YmL7hj2PidqrmuFGC
Xb0wiBgWVXcCGulQA/LvwTcHN2TAaCj/0C8XSbWRyJI2U+RzsMv/0JnLCuyfQG5rBK3msjRv37hm
InA4D8SsjqNBJ2lQLhb7hpmVJCiMIoxqCurIJ6aeVry3vJ/7VfbohMxYYxV89qQW3OqE1FC+MR0u
5yFInpjMCtKJ5TPAt/lYCBh0nL08rCBeqXDBTsNgUQ8WQgv6KPJVzJRWIIoVmQpnL/DurDduPk0W
4mS3rN8QiyPokA61Ct4MffoJGIKaM2f2AdAx4kffsVW8OmsbBvF90GuC/k5ZyEY9aSkBMVN3mP3N
Tb2IzWHFpCP6qGEcWU7dDBCKe64RL1bX8hlrtZmtESipJDRiDNupgCR4zJZbHDwmRKmkAoqI4ZF8
d9Q4Cx9qMgsdORCi9XOSNRpARMkxy5e1LTe38RhSbu5bYf3h/IhEeK3VnAEOCT/flDe6QRxjby9T
TKNhyIaOPVx+o/dqIZO+JwUqMxA76Z61MqoiBiv+30oE/Q1gZfjvfRMZn7RQgdskXuJLVpS/Xztj
9/ZfFnQM0s/dNkkuRMOa1+0N6WF3zwUJjJv/4juAYGMEiiFz6VZ2IH1gU1tJ3kcWjPlju+yABzI5
tVtLDmvKVV45dAjWeCK7TcKzAhJsB7Rba82ZPJq2zmEh1bEad1CUKPTUHzKfm+Nn7tecDV3ChH0o
gToha4bVHW1Qotv+TCJRRempZLkFCikrWJvXsf41TiHA9BOoieDsu1Y3KZCZzs1YXIf2cREx4ncM
HHWpEUnEb3Ryfx1Seq5baz+uyQh8T2xiKYUTJq+cw6N9ma67T5PLjmMhXW4sOI/pjtVFlXlo9jHX
5CD6wi+O3cgPhQF/qkDljt0f0hQ/Yugyb5Md+kgYpVcfzBeJebz38KJWVZZ0C/bPE37vrG4BHdvr
YXKHC0/jf9F7k5qOTilV3EBbnEWd4UshRyKQIP1+PdzrRYjxb2rTJxaxfxelwMPnVZyr7adE03lB
K9SZ2r2vIgM8Mf1oqVRy8ZpxGX44RPvXZMW+yfuYYlkzHMb+BCWLuvicwwkq/eRQVbL14LM0har9
rW8rRn8ZnxpSGr8h8GWv7dVsJ4D2bBK2Gw4k1Kg0zKs2hyestd+hku3rWWJhh22Oo4HE2513ddDQ
JSrKWU8ggTnunQh2K/cksotGDlsalUVgj5cd7PfXBt0T42QD/DYpz6rxmpQTXbhUpIEO0tGPIXzc
co5+JZ5oEzakRC74cdKmAikp26VhGkT1flGSYbevLmM/JDVCWHw+/w7PHdWz2ldHSbFnss+DsSL8
8ehveVRQAWkt7cRhRYMMXBNXWN1UA9vE/PLRWVG3RxKacaVE9Hi0JJ7CgvZvNV2Y0MZuXE0uTrml
N4CRyLY8rzFth76Aj6YkG5bw8SybYL8NZ/1+Xf/pY9HLKa7jwgIbx4pKn2xfM9m/7vqbELNpDBYh
haJIe07+q07ZPD9KO98uFEHXOuQOtaQiJpXI/LX9Y6U0BzcKc2eG25RP2+LYzVJjJ2jcYyQBhIKT
oStXqaZ/h4T0T7vaXPinWoqgRHWkMZtJT4Cg5ORSolnxfUvPADGx1PXkU5MYU2CcmsOYZXErb9Xl
uwrY/aWH+/CiV5v/u4WunJ7jvFQ6tJypUNNNCpShL2whT5Jl6UNOq3utN8TRq8sbcjSl7IHYRxdH
gp3I2FkPEVhsL22wSjM4Lo58hyOqst4rgRsbcDS77gnoCniIC/MUSrWZtMyrg2hqdR2LZL8l7AAk
UM7UAaBEvuxqP7TJ5YwTY8yUP9j+vx0SPrv1QpU3f4drtkvt1hxFL/2Jn06o55K7UBt+OSa2WEUd
z2UgLVCsdkizZrB89WWCxmKGQxqRLCVE3klEmjBf1CFMXXsDTAoRW2KAdVF1uMxKwQ5Sdc3rirOo
MaMONxxjO6ef/d1ldT95ZWKJ6lTTjUApcSrEpMiu5zEMgdYM8y6OCLMDvu5R5gq8mgWJ0ME/hYTt
HkscT0xZWh1L5PgekdxZ4iLYFjpdvgUxIROGkzwXckhLFBC6j9BJnehzkX0lr6Vh5Txw1TxeMUFo
eeY3lNP4YF0pxuyQO3sVQNIVcFK6tH+JiJKGo0+2Q6CzGE02j5vdWnFRQXuP2jTmuS0jX8PYlReS
LcDUZyOTnyBNrbPqS5xxi1B5KMa5yD2a36HGl60ipQqh1BttRLxDwzZUmMKwW/0GMbf9rtwWX0ej
0fnyVptr/jt112tHlc9cnSMq9BJtZVjRowfAIFuYk8588FPPjIXHd3vFRIMR8B/zcfMJOZRu7e1Z
LvEDblmTEeCLlEWlGr2qWhlPIb1xwPCKphJ+JOFJWSNvZKvJUOuB0dnO1wWHMkPUHuYmlO3XUcHN
G2pljzJJYZHatNk+w08PYvMP7MFcYpzZGJb9N+LBVDFJFKw+pCnhDuTgenY74xD/YyPbGy/VGcMI
jzmI1pg1sCDncS4xg86c6ymzamumRKHiQ+tmQ1umUCnze9zADdYxbuhIUC9HjyztzpeAbtpp38Iq
VKAfHtjSLuMU77HLG0bnjORxryerNpmr9crckVCrBYlEde3gbTwOM0OzJwU0IoAKbabeKGbdENJS
Iz1/+i8egqaGiIEa0kWlL0pKbrYCIe8+xtYm41Vy/mUtg7GHx6mcg1+haE223E5k1yPkQ3uw0Dn0
jFtkk1dzPpiHo9fTUcPvafF/BpeUE9m0m/g7wBD3FHTXA19WgSMTg9n1bU5z1MzofaPdanz1WhTL
sMUM0pI+59e1t7WQrSrMzO+K0ssaWDqVm/bw10RRktC4zbFAoZNtfjCNMjfnKvBoJ/rqkiG0fRBq
876lnl3bmv7/n+UBSqnkjqdSPKoSWMZWJDu6m6xzLv/kDw1f1nS+pOgrrrfYHzdtRJCMNsZuCz1U
lP3hQ7jmiOX+48yiQElIvhaOea2BfMtLEbMpLgNoLBqOBh9bEkw4UEVonkRA3tr288ZVNPJKoTSH
sPdlPly0orxscYyDK3YQsEywcznsr6rhFNLRn+Nr+KCCVKSR0IZnvz7386vCJeAZoL98rrwZwBOT
8FZJWDAXp6BqPYLu71bi0yWbs++KUorA6JIJ40HjfVj9kkPkMeiMc9P1kUZ8n2Acm4N9LW42FTxB
RBv5B9JoQAlfgn6O/OvkoRYXXYCBgKhgnzMfOvEsgLZGg2d4rjJzNasc4+UnD/hEXYR8599Dtbg4
FsVmw3+LweWE1V0qdcFM9pL0LYO4rJyVBLbc0DdMkjZBq3/5ONmcca/FarkL7XqjEzs9iWTJPq+J
l0Qcfy7SDMUFbVP2i9XoCB2Eins0KkGQEl0c/r7rpRxkmJraeFG5lKQhX5eWG3wxg+ZdbjEP4LYG
QRS5j3GC8kOXB0mYum+kGGDkQGqMBzO7pf5ABuIgJzWU+O1vAw8DINvtiTUKafuHLSocS4y/SQg1
VvbczeSaDgz+W4cSC5sAl52Mv471DotnMEAfeJg/99JOPPy5PHROe8mCvrYozuc4Z/o9YIrFvRpL
2Gw+yNs6u5wMNo7N+jjEnK4KHGMdSHceHSJjK5N6DK6gltI0PPswn8cySKgHQdRvcKK/htALn5zZ
/evsA0Nqj6zzS+Wr3uEgjbOXOxuJxRlInP558kRIlTLDDDiUyczrtsAkoXPgS1OGkhH3gSe4er+S
CckDqT1X/lqIQZlmhMnqbcfaUZ4AsVtDG7Jb3UogGWzMK99FZp40s23Fu5lL1zAYFj2cllft/OY4
YLNtNrEc5JnfjhzyYwOeecIeCIzrX+J1wUUf5EpDmGZO3X08GQkwzbD1q//0eY+W1rymfSZNxJh9
eLNJepbEmKY+ym2Svj7aKkMCbYxKu8ZZNInIkoFYGUn80fjwdbdiGxbj1sdzHo1n/cUaSKujkFOK
Iry6kSMI53OtqXG+MD7RUTSSw/DtRoxjvhwpbLYrWTB7ht5mxaWn5psWgEPaJZAbdfMcxjAVn4T2
MN4lHbpPEBdzvUQ1HdH3sEwpagJHeG/zrCb0cuouTOpJDmQtOcwJ8rs06XItEkV7nf8HRQhRAcCf
Erp2sO4Ggpz4L4VNQLfDcUfHY9eJuH36eNwR/p4yttGc7FA34hAgdYj1Ar7zpHXTbfHKBVvdluJ2
+NRrtGMOp14SAHq9Wi9xcxAWQjyXDr1Rq5BXJJvaboosvK17YDvfA0ZZh1c+dynNV5QaothwdwDh
PWdjgGL61kfwx30GfaBlLQ4yKdiE9n2VoUYXx5a5JMKYUkhbDKF8bB/XJ32zb8FTPoG0h4sbrpDM
Rm1IhjgJvoTktZ+ES0sZeoemcQ2tMII9Vx0CS9M/UjQU7HIQKF3rqZxcF99YAPtcELyZcqCOmZOx
HU/814gTWiHWBe+yN28xBmhV6AzQPmFwFh8GXO6VnFBypndIAkcPkxyo5wQvW8GSm3GtAakaauSf
ICTLKU23XpQbw/DNB5NHx8BlWxcJWFpZA9PEbIv5N9xCQgPdy0azBHxemFtpyTwvFy8n0lgeGC8k
YMy/ous5uEkimDYNxeI1wqY3mSglIOmVAVgGwW4cXQ29NtLN7nhEdIaU54/mdVtYviG/kDqKghfc
+8tvV18R+I9dHHnaqDGR1NLT2WKarC6Qe6RNUz+YVOcUjYrsn+6Qumb6EFSZHt9sgDqRcKKgDzXt
L+MYDoh3H4kMh/rLkJo8wzoMtN2YAr22Qnq3ZNJYnDCVAew8VFlmUSMG+YhSDsVxJ911IIaoJTIs
tFJMmnY8ViHRZg9Bj+6ZAgkgxoGtSsNMR02Eeh3lDUgchbIMq325jaa9sf04fGmaOUeFIw1XTHzL
weMPeiw6vHXeaKoFOlU6CEsdgcSulQvZ/4d5NuIf0pi7nKbfs1++D7d/udQBcS7lhqruYif8TLOa
0gferdjaB5UdsX3lwm6vtp7h7bIDkDIohnbuJdnZ3uWTkHkhOQUKZxJGer2RgyaSti98RsDC3NBZ
qGh18sKq++9SocBdUEH7K/6nXSjUBJUQV/CPvpwtcl1xCx2iRUh1TLkh8DvkBC++bxnKWlPxC1tM
jtaxf+gj3S+3QiyDQ0JjjZwMnZlUt+wj9Ri7wus9p6TY54yGZlJPk5PMZK0CjeoFFfpnw2R5sLlz
0e9sps8RAYXQiTK8CMmrxEOzGZKQKG7IKbWAW1TF8PWon/H0px99qFtX8eBeOnRrkCj2S8hklZvy
b48kvxUNwPqX35hlAWafpFelQXA/ArjKz1cx2/1ivfRRO/PRYvjy5Y+RuAh6Tr4QktDLxvJl+ew/
SykFwNEJrh+N8Lf4oJHZe0gtYwaUYxfSlCnOPUuYD2hoVAZ6g4vNWmR0X4VyzhrrsKiRow8EZbkz
bizAE8cIG8MGwFPqNoALc0qXcdmP5TLvOaktBAz6yeQxSVjRuMxQlQU5LQ/k7XEFXwEbt5sC2ulL
guVsKVnEdZ87jvAJJTHVUbX9xHgRDfNFiB1SHfJlDamyH9NF7CSk6fnFRmtoHjZSyuXt4d9R6cn7
0eBfPBADhyK1th2nGxhGV+20ZjyJAEki2NfGHPWV+JEGPA+N1BCAeiP+8oFYoJOy15Wo5fZjr0nw
CmDowrKKLofY3DcTuFrScfX6414Lv5iIz2gMH28okc+JuPZ1kwu+sgEHOSpNwgah9X1P/G2lx9S0
tFCf/VKtARVAIEXyNeJajyllEnF0TqvfscScSlSUnrZ7EJ9XNPewmbn2EEXdYcrySXrfDFxhQ7a+
5Sm42Vqidq6Z6hWSdIWITHDWFs9bmP6f+BzVjK3ZkA1C6DY01TPUGZAAk8sEL0kAEynV6wdAQL+8
OxkkFBEN1HrVnJCySJ7HCHjqMKo/uaTUtmR9lSc/8HW8Gj3ymJdDSqVSeO9XIGu4ytD0BZyG0Bzr
TUrG0IX4ozYbvUQjOJZ1/nnAEqxMLd5u00MAbGmMktkzB0PZsMbQvmI0PjEWrE/lVlsqbqOOplrV
j3eN20jT2ncFjidZZyGgConvSBghrSOvqOGa5gfuv480e4y0bh+ZrZQE4K+qF8LBX+7Sds8tJZCz
Sw7O7WG+TmV6/oA2beUT+HrpDs9fLUi2Ryvr1WDcNJGbuZsQfDB7Z6RpHy+Sqh8ds/U6P+cIT90b
Den8ZuAmLWIf1IZ1Lt9ABZRVNYRErymCsUs9uhtCmPMjwlZQisZ6MvBijEZMyh5xdtNVKvKuZKMV
UbsYivkf2KgIzVIPh5UKuiHg1cO/hjKXoV8Z7Br8ZoMQpcJ0o56ens+lLy0DM7F+M+bB6UCb5e6Y
leBE+7ofLO/8XxLp536sVzap0nsufoMk9uFE6ouq7WYWxzBUxy6zvz78WI2hgY2tATPfF4hVdr8u
pFsM0oLF/ElY+3O8DJIksLhEm4ekpV38Uwh/KR2R1rHe6nWdalNbYilJU4dzoXlSTRbuNXHhALIc
R+vNj7bxn0MYxeODpDdEW/6/0sM2deTvf6Jamg0/kkYiIn9Hei60O1sZGloMFl/Q9feoQ3yF+P8Z
4gVhugYMqS1rpom45tXn9jgo2IHdv+CLtW67k8VE9ZqAj77h/zHjkLA4lyaIeLfAYhGpfODH+a0n
F/MXp9HlVnQknOuaoYtLM79+GQPNYmrUSc0Dtw7u/JXm4K6lmth7uTEWJ9K8G8RpZLK5yKp+Ct3n
KnE6mhreVAX/Xuvn0C7RWPvMFDyXugtECaKGe9J2g1GtXRIGHWGdRiiaL/85RFCvOZu15jpEe/jM
KnMRSNJwi2B4pl4tQifJaBg9PsrCtPbH/bmKdWUzd5kyWYmZP/3CIJIr/Ohcew9DOlzt98UYAOzp
LexLcuBuG9e0ugHDeEUEfESilk1tIgdPzinquPo3ay+sc4r1xOrudCNzP1L8ISE/HS3B8B18yB59
lbDRsjwhNOqdFMqfeM3XoEkfquu2WwIkzXQ2gLQdBvtf7Jg8wKrJD40TAWO633hYjFXrFO48m4Uk
LRCmcz6q4Q2/6iE03ITnKkX+qALBLuTfRVKHmFr1VAVi+QrQQwumxmaPIEaVKcEBzkx5RDoADsuF
k9NTA3HWEBISEIUgvByXsCvEvksHe1cRWFIQDttxwoKJRumLgp4LfU8MCxTQUG0H+EGCjiBI3l7T
Wh9xnE5xLvIbcPAe/RWchsHBpGSN3+szb0RT6HJLyC/9zvouTZUpDf4x+UZ68qrkyTN7uoPFHD1e
vMs/cd8oIDVJVBxdzi0qQ7AxPvHxu8s/oVklJ6ayuQvzIVUdyB/Ihmot+ZcdEYXUXu/+sI7ACLOb
JR89xZ3j1RedyLJW/xdVFFkpuTizM4KtoaBG7fyp2H89F8/amKw2pd3pcNPVvzMR8x/6PKJ378cy
80jEG9hUkIgFOQhLEyaAWjuinwl0hrxH9t0zC8Zn/Ee/lLZ5VnDINtQdV+OV4tlDoAi3lRUIpLUZ
rDwQueVpjQGu8gEt0aDcK+lwyRwojQS/brcrk8I4iXuLzB9A8DFKvOLAV1vqBFAGzSup18pqVRx/
XhMPJEP8XdJGarvc8XNb5pcDr1SZy5eLcbhZ9dbW2ZfxCWAW0u1DbNTXY9b7fU6bTPXjGZd9AAGl
z6GI/ykvozg4dZ4LpA5NKMeTBjhlyccbD4AHPnRsstgGNi7Sq13Ck1hUmSICAkldAwArJk6G7AFw
fJwLZbym9Eh1IhPAHPh51vj+dwufq1E6Lej2waG5vfftpc0lXwXVn3ZRKNkkcjLlzza9BJ7W4ilt
GbgdtIaFb22DV3hLcdoAq5NYranj6yseMkQCiGRzSdtJQCR6KhIdYaf2VUoFTwVHc/paJOQ4PHh0
qJy5AZQGJwJh8dPNNmBcgkCzxNDIJB88TMG52cqQwHE08WF+sL8Kt/rAhpCdrpPSBnzylWRPAwo3
brAhZASFU72ptqHcEjXFXpCrath99pi6PDXKRJKRrLypiNGGLteqF+d9fyLFtaooXuXMndgZr8SB
TZcezY7pd6sGjjnDI3ojPVROpGgjtoJtwHTrkOhg0+jfcFZh+LwbynZhMGa6P97e3yya2J8C04cK
bCjrexJOyjaem1lGj42q2gJjcOH3/f5G16Msg/SecEKAfIiQNgbaKILqhaWZkUn7Im4pODhRxhzY
GjpLRh3nvFm9D4YV8D6oq7dZtEFStc4dxv4XfxzOU85NtAXvqyT9/390fo8MYAZt1qavb7cLxaTe
OLYZ00AvHGBb7KT4sTeDTgOOouPi0CNNSEVMVEEosOcDgE3LrMmZqvyqx2cud/ZidvXoEvhmRyqz
5iNVu031sqIqC6BWyd5HMS6TLITjAh99PuE0Cibx8rAP4RioIbP1w/Ps6JXoUpFNADKst2Wb3Pib
c0qHqsBFbhTOuU7BCKliCIbWTT0IJhHkqpvChn/DDJKTEDOXeMofX7s4nz0ZD6GQJHMNZVkIMrZ8
7ROSbtVqHM0qqDAqnJqfgYiumuWWx2x+VuXjN1B+Q3/MC6MzsItLc/Fd5+QMoX1qigg5Ci0L0o/M
NMIDsBJ9HdnNxFb1DvltVuytjWI2mh0UHMRYtBKxSNToFYMyNWX10FArkjrwdYdy0DfzRK69YIiE
oR66nTM4nZElOMQwMVa0YRSqseR9wc55sdFXmp7rkxuh/RceXeM5ylwnFghRqlCGuktKS7dQAPg1
aFZ8MUituoayiLbaTsLoV7sjU0DWG0j9ElvTuczSMTRBpFhTlXxA5PYYE0shoVuY5EjZUskTpPkB
CFpRbLEC/km1sxGcmJ1SHb8yimaJo9QFMpnPqPGXYVFKzDbaO0u8htzgBfEX9f0m2nIw7pwcizOd
MGI546pwyE7bn8dddpz8apsJV5ndpWH0ns3jM/oWNZ8Rj6V3cpxGc/2DGGVT2SxVtkaTXkgOz0mc
luX2rpnIPjOdT327SV/9cs6vOUgoZ7xIyzTuo1La4hELlL1LfDhYv9AQjL87L2bvSovWsD8gm4dD
nfNVUdIiVq06C1PVwdQKcOazFogYttpk75vNdI3zZEcO6oc0Ch7K0wF4GKmMWLlX5B894PJ/p7C8
TVpoQlmm7zCoPpjec4qIkzkZtjyT+PiEc1LjfFNlSXjz26OYbF4JKB/8FqJO3e1NtovUxAJ7t7jC
An45PMkjZS/zd044Q+GMHj1VHT14f5i09kKScXJtxLb32obRas7T4h+3Nysdi9pJ9f2jEOO3bWqY
jeTnML0jetPPrNGxslxklqwb+mFrQJiGvbQE8cQS3lAlqGeV23CqXlHN4EbLr7PY5bcd6RC0P9rg
8nfEEsyx1LWYe7SbFwoxKbQ1UIYZcSajOxeRaRs0Wbru8a+YTcwX2zluN66MobUpe4Xk49FQ2s3f
Nc3RfxxYAhln7DN5Xgw/1a+Ti3/e5Vah6MBma9xm68gVYc3c1mZyPEaVuQ2GAvXjAjp9p95JuXnf
8VdfcRTFF/d2NwRqziwgD9ZwlXZn0PasALKpV259A5Rx+y9c3wIlPNf+QImpK7zje0tt05PuhofU
qj/yy8dfLQGr3QL+a7sOYDoueomjrwoUszbKfmu18AE220tCQruUYZmogI+I/GCDNlUy/lbIxcvq
4pWyQCJeyG7pb+z5aoX63nk5C955v8YxE2aakQKBV6RF1X842JxmCytRk3BFr4ByFAaWETF6qij+
a1XPnxUzNPRTXPlmk2X3rFW1pvQp4qCY8/LMq511inh7w/sM6O64rXQe6Ij6M9rTTWw7lzXYXlOr
J6sYOh3u/uXxHrX8zeXhUj76wG0KDEaGftXE5FzXzQibTBcdN6iZmfDLlb56w51xSamODZ1BBTD9
MLaGULd2ZBBPKhexuAqcFlrTDQbARN+gbrK4L2800zAp/oHTdDqkAijqydqyGi/4wKQcudlpr4kN
NSU+E/2ttBI73kphquub90wklMlKReufFmLG/hm4jkvodiCqzhmreGbHSSRcrLPIMGgf6+r23dig
9ybjq2HaMGa+FkoU1RSt0SwjaeAJKjybwWzx0oAassf0ixssGzHv/vjbIc9OXSVM7yL2bbvy9CZM
t49ImNk326TqmtffOE+rB0Ooi+1QH5z0+ED61U4TT1mvccvN1X4J6psmLOqXQ19rGm+KWlUcjfNa
5V9aOuyyImpp7ejaDMuYQm7rXgNtOXb1BViftL+8pwmfp21ahFJ70zCZFRwnHHl0a/1GiIJnJlpJ
2kcEXishEvV+zx+Q562TETljl13WyJSlHx3BvZN9JDmgm2IZXORHRELorHHRehvr9yKPZsjwizDc
000DRwEToQh1p6Mxtmpmgr5xIYQ7pT2I/TLYlzU3vRlkYOC0AexuZ+b3FpOz68grLb+VvEqx8xii
OM8T97L9U6OhY4U/OYAQcWiQ986cueT5x8QzO9s6uQLRrVh1ZvchfJNNdpmmN+FwLFs4FZYsgCVl
Zy6pPd02BkMa6Lp1h3nb2CE7qeLv9GeSM2UD2DTMAgpXd8CG66xhQJnOzDGDvsQUzYSa+6JSGFrx
uOwtLTVqYUc6w/Q7Ogr7qSWq+/1YnKV9Oet66zrDcBQ+2kG9kxegqWSslDlbdWmhpPYTEulp45kR
jDgUGMjmTwTh1DeTnU3oMhu1RcbcqzE0lA8WMhw01s4z005tCBoLgzYsODVhYNa/0b/5BBHl2j/J
EWMwNdxf9kWIuLLgIiFkbf46VAebQyA957rJ4M2+A1kSWUUwYuaxNnU+mWl4C2TKXINt3AbjX9UF
d/GZQF27H2zFEfyzZGD74T/u6zrWoOKPpSs4skFwYouqka6349bsCxNB6x5n66jICSgyqGTvvH9U
Wq2MjOGr9AafbsjbC9RNkOGGK3ENzQRE/VU3iFBk+d4kzNO8qR4Tgr1yDoWJbevhpAB5UmOwJYFH
piafF4ciDRSxCNrBDMaNeVEC7GAmE2s/F1YLgUfZuxRiOQna/zn/MMqBJjRb2fT8SxSyzqX3seiu
ji+0sboZPoU+uMDrbDSaq2r0MWYLEaAOXaDHZDtAUOSwVvwzouRt/zvCtFU5Xd5zHd2tBZ8XAj8P
tueLWDgmPxqd6pGkFWtuVMW/uipyOxhCDhUWzNyn1O6jeEqBx+x7K7g07V/3a6AbwcWB9YMSXbzi
tXXAZkKjfxVHKwC5T8TnmoU8q39Jc4ulv8Sqy5aqUMsruaDDRNxxdwZjGcYTFAwyxP+EIldXomin
hymNm9isyuFkZaLOmwqyoZqCsn+9e8e5A1OB3qoGkoMZ00sX4JVujbsMldZGFqcIyVeYKpwbC+MR
pm+SdaGmosKHbyrFRAtlojffGKY1ypRZhUNPgN+NEJdv1aoQcSfYRiAH9V/11PPJn/2qpBqwILY5
LoTRFMqPgV31KbxbyeiRRIeI+kFjwte7cBhJcTcmRId1V0Ez6PkRSprsw0eR2Lcwy017c40PXP0F
jJ0aIj5Qs0nJka5pJCUybfdHsUoMlp8iI7aKX/fB/OunqcauJHHH/keS6Iz4YsR2BKuZbZ7I+J6O
HrTVD0wxVvxklFPKRxiTH+pIMt3rn4eTypUimMtbVcXI8FllNVdQyIBcywE7iYXttxDqHlDa1NyM
kEgXU9d9ZfoPuXo79XpS8HRF5iJsc6n8Y5MupoRruRt7BM8W1wFX1KDMNJXx6hbXpVcJlst3SQWF
HcBjeoDugPBRvXIUDp/95c9n8FbBsHRRMOO/QDvy5EyTT5zY4c7ydL/Db8y9i/JHryVHAu2PtDdS
aCbcQLE0Xg6Zqn1Om7D0h0wn1huaITqXOGHA/YYtUtgvnafbciVUFwTI26aomIdsgxcFhpUBXZf5
2mCXsmYxJUz/EFsPmyH/hL0eff0I8fSHJRF3i/sYWyhYWyGP3UqP+hBoS7pRRKHmoDPDk/GQ2Jg1
GCMWf5g58eVTFmjT872favUwMFYujhfd24e9yCqIbOBUn3rjZ0OPSU8wIw0RcNnT6GX5yA+F/90b
WlcU9D0aYHRIyLMBj4zwBj5S1Eiz7eHSir6Ywdrs4zcu2/ni39JaY6niisUh9Om7ci7TOMKVYy4J
2Ng4uU5STwnFFl5bII/MX63po5iVArbKVsLda+FnxzhLbgX/1tk70Tl9kNrXXofywI3CkR4xG0kC
7E9UqOkLScxsPmLuxJE+En9bt0T9NqKbFUNHPO9+/vFlRs6ods2x0scSP5RmzS9NGzVaAdWHlPVg
SdM0DQiZTyIrurOvnCDjWydEKyMQT/9j0evIxh2Z6mtfBrRQ68wWbFzwkQiEiGTYNZpjJwQmykLD
YrrMciDOYIC3ZkG0ixDBXvJcv1trYaFqpBSGspfUYZKsQ1Vw/KWM41eCS3HEr+LAnC7nwvtAWnZn
XJYuCVx5c35j4gtXoJus5rhEuf5dweDkHtpk2zp3MHFO4oU69mhQ5W7jZBYh0Ejb8MJWrOiBquez
U30lzmw3Rw3IXrddfsJEebQf4e0JICk+pSx6mas2YJekSZV/dNHxNTRjRs1pMh76s4ud2MCLMf58
rT/kOmX5Ep3g+ufCnbL4LibMg5ra6OyUNoYSgtQlvzLyfokjL3k3UgShacNPlrHtUONWTc7C78nE
Hm72aRy1J40ovrSKHdoDTRh+Ugn+Zfs5siWGiJLaXAzq7HgIebyufQkPbU92Di2ecZ97b1qZBaeb
8HhJsH46g3YQwok2aaIAs/9w40oDdIHGCM9aok8u3U+IiuYl/8zWPPytm2TUQL3tppYfkB+Qwf+A
sN0U4fKM1ixVq58sZq2LMQjqTRSSnwJksuVXpjfd05ATR9RXUoCwGic18rx6Nl8dmCWeK4LwL5zi
oLsi9dW0AO5od3WPuJvkUluCO/G1cK8UUXhWTHv5ZtfOTUw0sypqEt3+0pRR+PhKa/QFR48Dvbjy
S2eBxJN2nisrC5OWC5KhywOndQbTKArMYkJATo2/OEd7Z0+Qmaef0+5fU+4MPSS+nLqZuv3/w6u1
PGPrSKWcBhQR6gIyQt+81w+83PAL/iSXKWiQ0uG0nMYhnlVjenByiLu5iEtWS1eHBg16lDin3alI
NyV0PvnpiwsKMCR4lS2PJBM5lpAt4ws96rWXftgRLqUc7uUdxGa8FD/J1gzrqwnj3Wq7GrtmDAP6
mXLAVqvUN6sitp19TP2cGwo5KSvzO2b21bVvXKtfEYzbQ+2XejSXH7imbNg2virybKyfaspCkrOA
NTiuA1U1jxbyLDQAwDwfYbPgfINs+8d3L5D7r0NfL6O75NoxzpjzLx8tyZ9lk7YHOH5206+/FdFi
Wa0Z6oGV8m8vWTDNAo+Q70EEkqAgxKwD5qrD3yUZS7K9Foe+HHhFXFxcsZXrQCVren6cGO/bo96q
7lUCZSm+CcuHSPi6yExqS85Ol/6mNtioV9mxqJ++MJ1lNqD0AAIEhsNeHzh10qD6w1IsAVuw/QvE
EHvH9dH0J/jQ62nSpA6cfcFZ1YR9QgTDgEDlZESqfuDO25BWmd+XviTc8f0CAUqntwhulnyMqFfI
kDihtUZv3vpAhtNkiqzH99ibj+X5x88HJKLnHK35bmXeniBM4xF6jk1lluv80TpdkyFhzDc5DPJL
sYuNxPoePCOkozFtx1vW0W32B7cJrbdxxb3w6TS9L0qoaAxAKeSy0YlUUCaAvSOy3GBkQHWAO8V6
Xcg2gf+VJrGtrWoj2pSyIzIOrN2VLMVUFlGeEDqPqgUGdbxdNaa/WO46fgLHSdxiM2hsYvuLr+Qk
9o2oFbTQdX76XMjZUJg2j3WfKSS8B9Nhe0icS/1rw3nSp+6zSHLajLqmUg5q8stZHJeAT2AA88N2
xQLVWsoT5a6xVHq8Hj3JHALaFIdfdX1+ev+rElX0EEIU9TG50XnEeu41cWoJHblcwM6Bi9qPsNCm
gETJjsITmMmwECDdYwviWnQd7S2ow59K8tBF3BpAj6akXFipHnkIS+sgV4AkplNh0Nhzl1A/DxX8
71oFbzabWx1TdzDRlz9n4BadP/ou+NL7Nqunq1FvjgfXKf3kIJR2adFjnxc3kJ/E+kaJj83Hkdb/
gV/KuHlbqS2CV6+wfLeUqIqL30sM46vEpxVAqPFNQ+gMiTiaa08+yl2uxixQk8Pl4FO5qHqUIZbl
Vuqf/Fa/uK6oi+kuzIrfCvUyFZJ/YfjVaplJyQgeuvTkuKwuPin+OGDvRcdgbFEt9pVpDx5xpiXB
L33zRke5xnBikntdipf0GgKx847gTV9osRu7oS5sSaytrgYoUSjM/eLpd+01QNemkEIbM92S/RYb
JVPFq5fe/MKT5IrkYZkIxYlCst4tODCOFaXUMkC3XmleC99kLSmSD917ROEVxTSa95xx9spQVuz6
l9j/UeQ6ENqj9nh1HESV9dyqR16D0lIbX3jz7W6gLj9xlFI4qX03/OmXNdic7n28QSjU+gmXT4zn
JeuMLo+Xq5YnUwB2zr85YyaCUVxdvViE6oLcHRIDejapkjP0q01f4/HqSatKgy8CgChLTvchgmvr
a9wo0miRrDyKg/E9YwEumMDd931OfAuCAe3/bBl/YKN0M+z6nMoAipP4zieN1QczzbX8sqMVWwmm
DVrKs45mCiRLKXGxUv4QqFoD0ug7tIuYn+MB1Q8sdiX1bNh+Czr6BgK6PjG6wKydeeo4m7ge79YO
U0aHHQSqlSMSRvEmbZ/JvyQbJK47whn0Iq9e/AZPiCrExgjWWipu7PGh+InxRMxfLlWMDFVcs90w
qoF2ChyNCNIpWERZlXbgQnIX7KwHtMt3jrt2dAykUi/zEeX3dfO7nDlJvYV3VSAId+WGJuGmBY8u
FdxBn7bGz0WkvEdHQ0tItiUwXZgrIgwDXqBK+NyDo84DkWtP98iFH4qMyspW76izY8Ikn+NWr0YO
efzrgqeDOaaQb0ajZFpQWOpdc0CYbCbQBWF1HQzrofF8g9DFx4WVdtVqMo7/QLAF/MX9OCh3PEdW
W/7JgwLKcxSMEzZyt03rXR2ie+iElzfdj5fVIJrhf3imtZdtVE8O8yC+f3aUwJVZc/Tziy1ZeCgw
ayKnBZ9AXRUSU91IyBCcOC1Nq/wDmc3ZCmgdNkzLFL/YLfiDmXNfrDQmBZ5GTswRW1jYhhtOTv7y
mz7bNOXO57f1nmfvr82n6FqK1iphhtseU+EHl7cIMWL9tpAATr7C/9tDqLJUDEBwyHufEbMvwHLR
IUbgtp4q647v7m2sK21qPNgX7wMp3/8q3K9cn5QcL02sMgEDj1iJm/5vavoEHSYmCXQ01MmemaGQ
6qaytgAIa6nPVIMcYkxrSUTajq5bQaXl9XDo3qFwR//EX9aIietJ6D40idTUq0SwoHKhUkLX8GTI
NGD7n1QfoaSU8U1bMMmrBs3+IUXoduPBaTAPK/AqC3z5T8Xn1nPadENIisq52ixkPctDYJ8qa9m2
RjuexwKmVxKGO49Wnug14EINNFTmibUK9CVoe6FJ75GQBhULRAAdQWGPKsdDqQPDEFZaEGsj25Vj
Da+nF1O2uw/oKcTSxJefOQpmDhW9e/eW1IB79MJo7BdE/BbbzGHmOV73Dg+4O9P4mi1ZV9lAM6Es
vOEF/aiC1Z52OpBmUXQg1C5nC7CtJCy8/QI1/gq8SyExKnWTE714az/C1oxfIsRW+fSWnMqFsyCr
5pnd2vkW7sd/O2VIM1n17JUpkng0ox+YhA/hX6ahHnZFOOSt/ZvLP9Nr5tsVjrjEjk8w65gCEZ+D
XtbCMSWJD1G2XxMTgjHDI+nMQo+BVrslYuR3gWESapCusIm4ngyL4OIxV++9h08IGhzONbNHVlx3
ZEnJyybM2f4D+m+VVYelOmU3jPyTwuzAyB75OMxtK8f9+G8fClQob6z8vx2PNJyKZqfYOqIzF0CY
9VjiA4o8dDTcOjqd0sujISbK6KCBOxpzsVdWudGe4pf2se9Dpamw8sIcgrEu1Z2oDXcWYxqzEYfD
WyoXAvBYbWMSkqJfVv68hGtDoteitPEgirTAQz4sUBUUj5LDLefUtRnxI/G98tcnoFptiZJRp1t0
33evibsXqzL1u6D7D5ucplYT66m4nvjEuqU8GD0RqNUJEf1wOF/aKyw4tBmBk0Ap4o6j48j0Hbhe
7jlrm5/QQ49NVucai67AyHywO/f3hV6/K6Gvh2/sQSVKO3PLNC+J4m2tFkZvFrfPo00pe+X3Zb79
bMqqLDeJW5WBYN5qZWwW8mQmim0Sa2NO5HbJbd2PAri87nwNUD/p/p4LrobFKC+DS5+kerd6NOxd
H8dr7IJTQWh1aFhR7x3pgqV0hIyTHoAiabIsuksph9zsohk06qTU5jL3zoAHOkwZaVvjirXkJCP3
8jWVh+4hS5ohrD8ZUGE1lz3lS/v+37yx0kSXg83+qcp69T/9WVuHHWTZaQblFLJTwhyItw9eyToE
uq3DHNRQCgH33vorF6rgnaU1pxZKQlXe37t98BEWX9myzQHeMOle1XSpU9gc2wD0QoXKZeP4j4Wj
sqz89gx8hAXjPeoQoVwhGuCFTsQ6PC3xqxU3NzmT/vRY69fgz26xeg8vM4cQMJ8Z8koTeqTsfKt3
F3uzEGWf53/s3Gzzu47aUTT2dd89Ovm+6+iPFb6XavotW8Wvd/EdEF0hjX+AV6JSWw+X4wrqk3NS
qJkq68zQROjvRHVzpbr8gnvZEIVQN2w3+RzUwFGZUlTTDUmFZi5qQZHAwREhvv3a9hG4bwCInhgi
EG9ScOaVxS5c+gE9zGD9KqCwm4GolNz1qslCK3c1d+9nRCmHOie/TOdZEQZhIChE8XhGZhRGJ0b/
/LX6dhh15XgTn7/BeCyP0BV/vVyshaRxWxwLrTptkxm7ZvRZia7DkZvGDnMmqS2puj8EGDfDw/73
OIqba868PZ1ErqGwrC8TxewUTH6yr0/XQX/jzCZ17pNTX8b96+HK3erdQXnLVfD2pubA79Cjvcqd
bxCgGjzqqwp/VieK65hjKSWTWYPm5ESE8jQ67ka4HYabqlkLQAU+YjKtiSVu8Y8h6YqPPluVMnqf
ZPJaFEqDyaFH144yGo6huc1t6lcQcvH4WZdfh1qct/3m8mO30y+iAdOvJinNHIg3mbD2ZRsi5HzY
tCiryEGoRPYZZDIu9h5Bycz1GSt+vfUEKtRfQaOeH17BbNFHbeRX+Ce5w2OkAY2bSYmS8roY70Hl
bwRhECzGd+G8mEsatQg4jvp2OypniF51slP55Vnoe/3IQxZrChTAGuORr6WRYUJdGY9T/LE02Tax
NuGxyt3EP+Kx2bTXqqPxz90pN1fe1CiNeum+gBibBthkTjVcB6bO6qukXrZT/vXUbHGKDVKs7jSF
RrXwzxXNzaFWHX3qbwUfxCcGvXZ7DCu5lO1VHglWw3QF9FDQ5hYzdvMp336c3GO7VFnQGyLKEWld
wtpDesqh2hUDwt019eLi6pUNoxwfl6PS92Ccyv9+AMRG+dM/mPuO0rnpWyH78sbREA1qtY1CjcgT
UztMMGMqO4ydfrVkMaej1JTvaeB0XeTVj7HwO3q58wbXUqjqRVyG9aJ4WHQiqSEKPEd39LfrZ2/m
o81klYWu2fE3RAqFvz0bdi+PE00VVDlS/qvP8AEVs1sB7WhkgfAJmrsNRV9RlKe+mabkW3S9bcgd
R3pe5DAkDqoFfHsKiY7x4O9D5OFS1Nsozv95NSRshB+COCZ+UQ1pOVq5icQ9cQKh0IbF0IIyVeIy
nHrYAPB1aa/UJ7FpYAZXRPZRI0ZTuczJX/x1ASxjUaId7ZL0XhuwmVUBnS6a/bXsAhjcvDCSv1Rv
Djde1xycSY0YAgj2UOpozZp6qaHQDxAg/PrhHHeolNDFw2DO/gKPCDPMs0YvBrVFi+uc852iRSc+
Lvh+CrLcTqQpIUj/qd8npbSu/5ucebDEkgHjm4mcSAbYv5+31eXeTQBVjBEFBwZDTKeVs7sSXVIQ
SBAYL0jPcdjsKWOICxUGsIchVgUrHPuKMn7Z+oJe2SkpghNzEfSsXi0w1M1g5YebvTkOMtaaC2N0
nCxKQIst2nMpizEboZdxhKYAyTb3ePuOXFqrIxMWhu/WSBRPhuHgPcRps3Mn726idicfwOMd7/T+
lYtNiODXspLxkGhmluvflos+/wvb7OvlBZ2ViMtDFsROEePK9PKaqEA8/wiiqZwtv4dHF10wmJCq
TOEmMIgcd2TOKpfv8fl1mIkkurvbUOY4bJU9Em+WZUto5r+4GGOUIAnGoUXhYRmHR9jilqkgEwUM
deyZMgvwXIBf9GL5ldCUY7pGNmbtWaD9E6SdeB+oKDlwg9oIMT+XbKrueH9V+wxWneTdG9jTkF1w
Oymfs+srnwr5v/Wr8/m9EgbqW3c4y/L9WKmdrCH+aFC/T0e3jwZdYIi+PT+FMeUINP1cgYIdLGoz
BfSTW12XkGFWEoWfQZ/swDXgCtJUxNDQ24eOrxLoAhWyyv9Har281sFYNwSZ88oGSfTZpVI63ONt
S6cMnNRevzcsWupNvKX1sjcXbzOiV4ZDZoZM8mlejSCd/eUVQD+mIGAtqEpW1cMVtnNT5MIgKAai
1vs0lSUUnWcjwguBQSl1+d4tTlJ37HyC5KksMs26K77dvmfe+yNfZP1NwnpOuJmORMu4Spsac8Kw
yZk24J2nW0fQe/wugslOfnACvdnreIdjp7NWfJ9uS+3TsvLnah5PPPo3kbqtEbkUKnrJ1WaesR0t
uG0t56Jarjz71Pw05IgoP+HO1AqKQ82VYbbZiyLQVLRkquNvIIIrBTaFwPrEt0kPf233WnCtQtbx
zmiot3RRoXuzqTM7gKXkPKtxPU236ngNP3ghc1utvs7RU2Va1OZDzM5aMD72BjsStG+yPSn6GmwS
x3NMrothUMb3wnM/0uXGJjc+b9qHW5pmpqq9ECCzG+KENfqVP2vxipWGUDKN/y2iKFiD9Lmvl6I2
ZunOlBel8vZWVFT5KsgklEF4FfvF/lykA9SH02oAsC3ghNbbjw6GJRTPGms4fKmwk+T96gqi/Tfc
whDnwfgblLAyx5JRCO1am5pQRNr5NT4LN1bCgesFgdl0rJ0h4ulx2J5OsAUyTQ12prZ3cvs+QZYS
uyIral1YqoGHkrFH9vERr+9XsFzUvSe2/Q76DPqG8xTPMsXtJJVOlwBFN4vYzU/s8b0zt9RXKetx
Ap4xvDAX+iQYE2ytgjLszdpLTedKDdksiqYZs+0wtrba6CPfDu5nF6cfcbzxjc5rtEtqV28N4Dda
SKQ0zZmBu8tOjG9qGviqMzfZUmpTsHQl3IxKstbD7keTPZWkpDRCYGtjflTNWGLFfa8TqDQSJ8Sg
NEB4WkixhDTfJ+WqTGziMrCV4EwU0ffL7mAMH7unSQOKPlqy9rrIDKUQQX4L/WsS28q7QsLw0sgo
8C94g91F1v+mqLnxtYqYZZEw8HE0VCwt7HM1Gb77Oft0+M86HRm6L3K6JrxcZGN8QmGuSHw1cKVs
EWLGDHQh652qy64/EWV5OO9N2tzVr9bf9vABDAKoHOx7l/fzUrrKlTKBZD77GBkN2IE1tT7imEvH
rfjTgxNZh7rM2o4qfSBjCfDZzH/5N6SY/Yt9MwRgpJYrXeelXPYEKgKqUAogYki3eIumLK7bnkWm
HCpq2ExmldmWusfxuQZ9BwdbKTleDZvy3Ayjc+qHdUA4A5TpVSs3g+8yAQW7trHgLi1MLVyiJxWO
xDdJ/HnjaDeK3JQ+Q2odIs43a6Fink3p42WauPIAuUU5PmQCCAgMd6DGUBMOPK5TtnP2RUTk4nTA
0rJwEjU1f5mcWsmblKrbvGBbcttO4gRYe3SQL1FRZ4n1qB+um6+pu2XIyK2E6MMQFlYtXnYBCegP
Dmh+aR4hEb0a+gv9/bIZTzwe0ID75upBZzHJntkJU2ATQ+7NahBsjnsIVmLpwdF0MOBLUJLvsXzq
KRrVp4lglHBwbm3a5s4Hqdg4T/zj4CTeAJGDXxgujIFN5UKifnP+Ns//HGuI0VSyO+OoV0wFaxnS
fjyoEkWno82llhuSDob1p6RxCbO7U3ZM7Uw9AmmnNzxjdxjkCueXKVY3mm3pbuyz4siscUFXSC/n
FqfsCGqeABe0M51ZN6ipPDa/tBauC7rEnrDZrur7ebtxwOZ4ohA2xLorPZrehGo/jjeFcqUKKzbg
MQUiRFd8FKlh2KCTB9QicpxuhKefN+bLV8KHDP+Aw016y+Ul8BQsssCYQFxZ3rXtjcODR4y4Th06
6E4lu5VA/gspD3cFDKCIknVetScq4JnHs/TjXc3HW1uW2wiALdvciyHRCGKEw5rA49mGS8BGonsA
PNg8f2HD4mJUTZuacwR0yBdwBXRH1zefqLSbCW98Hsq6rupD4odKxTr3aKyXWlISgCbKZe26XVv4
6fxpBQ0Xegx/KKg2j8T/0dci9K/gVo0fCYE98clw1ocXLUxDAngZ44ko0dkyc+pnaTG6bT43Rle4
nU48c8BltP3dVLslSKjws5rPuacmaCUPWJY1H6rG6j9J2R8A5qBHa6Q+CRAG2xDoB1cbUFnuBqIt
2gtagQfjYJ2HAYgP2igaF3/AyrdXtMny+8Th5dzadpnMm48WVfM4sF5vvjvxcFpos4PvME0qeVLQ
Ney/b4WXUgGMSBlPqJ/824uf2bIGXGPaoQ3Wh83pGO0gZt4MnlAQrj2UVXjoglBlGT91JPW2Io0m
NOoqVfLlJ+nWMvhd14FeGoOyu+aG17Grldi8uZWwjqcMX0XaFlVMbozEQpn+swqgYJoELtnuFJWs
DR5kDBQ9EF6SoSd1XuIV6ma0JvjgUPSrDfj3DxF4Ou/b1yDX5BcIpbWHvmgAVXXHFUptI1SPLz95
bk46Ev01VvYYSKqgrxl8yJnrV/PCkbXvr8zfVH8X+oJHBbIO57SBlxZW4r4ty2qgImSq64OjkqUB
gifFHAea9fmNExqNSNLecl+cYXznDEbJrf6KMqnBQVR9VclM7L+gdJs60PqjTNTvPZ8G+0sUG/k0
pT/AWPASXNy/4X6kttMcOKIoUH/nz+5+Lu1uasSC4HgovQgD8KvrRqC0FvNxEn+N/AsYSl2KemHm
76Na5RZd5qEjeE7IVS9g7O65uNisjsgKlW6+gA6bQgHOq9heJNsWcYeccP3cc3posIKT0nMJQggT
WmMSMLaaoC3rDuWiZ+A8WuDQy/jHvsFKKZJpASvIBT6vMjuz3b4k1oNoqpmgEiixfr4ECChT/a+V
Q89ND+zZgci94oHdBgXmAxSFR52sKv3CPsrW9FWFtGcdJOxUxNvDG3+nolHYlXSrxJRoemNw4iJL
HbW/SkRF1x+Kce0yRTxPxT2vbTY1c7EyD2qxmNA0CAyt8DTRhkFTYWtx5Fok95I12I67m9Im4p9Q
J6PhFPdp4bEX3jDQ4ChDgm4Qq5JLAuLi6OvxFIska8+XK1JrGSW0lzyIXncwuqh7fGmajYBnR3dH
1bERS6JD8/cQSi8TPT1qn0PvyqFu+lo6KfgNfZx5l4dGy/6NxGG7Vn7Ll6UkGRoslQhSv6Vd1sO7
ubrNdpMEIeEzCb2/Sn/veJgnRiqpECzBi0W8XYW+XWEoah3hYd446ErRX+yutdMcz0N364oZfayH
PMsU1CHSRXXeNgOQuFWvabOHZAZ6HZg5biZmZ3dQf60NeNSO3DG/jBSNwULeLrQEsi2jNRcvy3A8
h/Ia7KO7HmoYZ886AhJtyuWGf9L+AnsQp5A7ibGFe4YezYJHMbN4HrEy8MJ1HGJVMv41GPuiWNx4
1sFLUalLK1M2MJMmTHaxswc5PpklMgwbgdQAgZ0Me8AnEaW8jSAeecz2W2LobEQp5NMjp2cc4hTW
42DhkOj80sFCOQj7N2Gwtibfnia0ByfABom0+eQ0PBDM5pcS7gXBdYVwYsKMDHtfDbDF/kx2e0/r
3oFrkoghovgtBEeIkAGYIfBzoab78cNi/5oyx6cn8Cl7ibuR2xNKFE9U86VoLFYidIeyJFrot/UA
59ZHtd/wDLa0Bp0qYtxtrkwUUGqwk9WKkmVSjCYjUDCqVmAZRTLI21dWaXRGnmrK7iWNE9KImjes
4d00tvouGNOWxzSTXefIAbQKqJKM6wvngck9Z9DdjM6uksPj0dY1CH9yQDwkBzbTnFrIQAcPcm1Y
XeJkJ5bzRFlJttDUZA3m7NmlfMpmCQjINGKwILqvbmZpAM5LGTN7ItP+tYWZHP0g5vRiYAVCYQTj
tH7R4/yrdxIzrnfotKes8x+D7iH2o4Uqyi7XLzZNqi+vo/bnOIkU9kQd4ccM2RO5udccSlnYtUwv
FymmXQHP89MtSanht7+RkB5Ig9XNxSyJSz/Gm8SNyn1oHF7rX1TUVXwDREYllX6JVMiN9d8A+4zO
5QAaZh5+dX4UGbxa+ICHvP8XjDiq1Gf05o9p07of/BUr4El+b4kHGJ7cEROOCIK3rBbNSVIo4/6K
hUt/0CM+iWCVPvcAhW6QxcF+aRLpUno5K5Y7LTdGqvw866KXq/Aj7cN3TzJKjJoNvrow66IZzgch
G2fVFuIb08Aee8o5V7/UHAovN0CPb9HJD7Am8nTLfgKS3rIbiK4JeizEV8UuuWKoZ9tDrOGyQz00
RhLJwR5bn2P7s/RSBhcIPcdlvdR5k3E67Xi0lyEiKYgEntmiviaLTlb7nYEGXr+zaZLWg+nJ/+oP
LW7t28z6odLtMhWFNkWusr5bzG18X0b2AeVnXcxsMXAuh0pq8Ysu9jMjj+GhirUDXWySajSCpQ6j
ERiPgOUsnMYOP/o5vKHgmIhfYCOgfUameol8NSwJRSNc7Si+1ZcedwbixvO80jiiomMfakOvgnLk
1+YW6oMBw6fzG9R1TNE+MMqfwIcIXFCZaw3nijQoNEaXSw/v5W8eS4m/cUJ91eqbfEm81H/zGBUu
TWlAwD5D1Ex711bbm7ymeuQm9PBiH4Y24mKox0k2+7FGDAGXuvL8ZUVSgcefh0WjXBOGCFs5kF3e
HlgMRl7TqJPvPKkUEJNKwoNJpDcQDmZW1ePpcFhdmeODughJrn7xGqbpbxr5hZGT6AfGoavzAmOY
zkO/xxUhCkgda/NvpqE0XJF5iYyrMfVEbsjNCxbs9MwRVmJHzOAQusWeyqDfDQ8ZZROHW4c9TtIe
g5fxzX8Gz2aXVNjmCxE/G6Z5E6B34iiaB8Qans2TLbmTMsASbXS7Es/1F9bgrubU8A66DnBJasRJ
ta6EPHl1JM3uGzMLTA7kOZIa4MK7uAHJP2H1OzhRVoa9iKdLQtEVc1ni520nrhAOsBLt87MSKlbD
oBA8eTwXtTyvqCI1fWJZ2f1AgWpD+WJhB8Dg3G/YEqTUsLicxpkqzn6H1Dv9/JtDRbpZ0M6S6hUK
t3sCwMb2URFFxRJiX+z+vjt6IFjfnCnjQPRvtmPUnZxDWDSVdNTdS42zBhOZkvVpdNk7OT8rpg3x
1s7zdKH8pcMPU64oLyoOmFHKrf71h40sqRtWgg3Qed/ZDmGhD8V4ztI2zSOEk9SrTHgw8UDn86Ki
kKnbaCC7RzZpjhc6mQocPBilm95ZnK2vmLDbHy4yzlPsOypLcapU3TCtS+faRLKdNAzm8Ne+4MtH
Wv4l+mqGx9YXfaZwq1gNegqpoPSRVlHuTf8oNn4cTd3+tS9ekDBz+zG/OOgWegrLpNf39mElZP2/
DOnvggxS8riizdZT4PObffuf0xnrH3tq+grXsAYBhFWsSDGtdLcZB6wAHyhiSSZUfVzKnTohL1K2
3uHBgezzfjulEM0r0wGneRr/lzRskZHrrxkrNfI5J2IDeZa2SZ9EoKRWIiPhzV9EBi++Yag2wZb+
bzU24HhKORF3D/eeJjVQ3dmrCW4FvT3WkjzaQTYHn1eOCls+kGby1Qv1OFVN9pDn3tc4YoSGNQBc
gBoja879Xn3GQrKtZaacCe21WEcKz1lucdd5DN/unF7RV21P9CD2F+2qFHOWOEUoCax6ipGZxom3
d8XxHbjwGitKkJv/4l+NYu6J2XX3lXeiIluFZnAQ/cv/tjRnUVxqOUHMdmGYfR/dyz6fIMvE51PM
t6+Hq60P8Im9cueWEj+VqyBWNeYnIXdWF2gx7cV5bHX+lhxO6eadaMzU7Ne0YYktPkF5wfvFHLn8
8ub+OfV+EBF2REiGMaBuUHGvmy+WDg7+xXBfypDRbB6DmoJSMwLtmJC46Ws7wErmnhAG+XK0TfgX
u9OQm5BJsmVmdvkiE1+Um1okoluwrsveeTOMrSPwZsEudZegrawTDJqgocly5Pk8Hzyp/cdxYdXj
mif+vS/pFYOLBmN/vqnVtyoqmdUuHiuoSkuDo4iyAHzzNzGHyOj2gO8nukmeZ1P/t5asQmnJVO35
8wjg6bTX49BY44cw9YzFYtdYZqpFKMGjmdk1ovCI3KxXqd3ISQlrQThuA6uQ0UPUhZzkpa4sv5QP
0Sc8MwsljOK6U4ZXLmdJ86x7vwxCoGD03wimeIp0l1jQ0MFpAeD1L3kOcbMOSJ89Y5nkGKTa5pgK
1KaqzYj+LNJmgK+I3m5xYiYzOfvNlIKyYj3qBGgWaTOxYlkSscFcl6uadlSjMjjEXJqQWM27A54l
PS1arv7XtsWdAaS/9XGbDjZISmXQORhnEySkNutGqZK61+/nB8L7qBDKEQLzno3jWUgDeQnP3bIs
USSleNffBioBMSknxUnSLMZauqW5N0EWdRwI6yjij5hO3lv+KnwxqL64h7PTr8CxkxNJa0i4Ff+A
79kBlIwx8DMpFMQS4TFEukGb+LKe/Bixy+lM5wDEK1nUMs9UgKCEXVpy34RE7IR44GbwEpdWtZSq
RHcI/a6EXdA3/zb9IDPTCwbJBc/Ao3UiPRqEbg6B6OyJQ2nfiE3h/f4vwLuV12uZkmdBne8VcLuA
KQ4rbJjflrdaPtL8G7bHm1IPUL4vfCFNIdi0cRxrfvj94Bqd+IxVnVMl+fW3y4miqUdNg1SgHkFH
0YVaS/FXPRHqvoNFt6ObNflRlUt2pK2dsUyKxMCxrsqNe4sLuZo8UWZNotpcamBlODYRmYYjxwdp
I5kIt93P77kPeTtjcoWN7eY3n7WTM15/wOROeSeY0GXlT1b+Qmue2ptff6lAINeCEU7k09a9QXIu
xM5idtk1HsPrgLDqqWhT7B+vTL5KNtHZY0tESgD65Jk1h2u6BYaOrKJ5pDdIkw5BiusWe7BgvakP
YX7UbxDcoNp9Mc0SHPia+gW1r4RB9Uba4P9qkDHimZjfr0+azxt2NcIidsqTq4WNwFWVVPNrnCW+
cVwxKSdppY1Fiz9vOay4z8+8K6ScTroDX2ZAhTpKwHJEyTDkLn7Vtfsphyt/+mPdvVEhpRmP0A9l
cu+F3cjPjv24F0kqHt63t1UaeNNOVF2mQVeWM4ZyaqcDnvxYpXD6q3d1eLVv13ujw4M+NuNj0FRX
1JlV6RXKxbI6xDjDJ9heCabguT6X14X6EbQN/fFruU2Gu/ZMJ2DHB2wwL35nWWoOUMPXavoThdLe
MgZN5T7YA2XgeBwAHCnzFrWQByTac2vqao31aCeXSKXoqC0eWHncrg3SXU3cuwSs82Qy1GanrCq0
PkIdi652T/CAH51PsrYJkad+bfp/xOe2REWvMt2QPWP7H4btd2GCAaMTXprvqlKAz5BXDr0d1X+w
Hb7dYWu5VrcIi8bPkcPm4mxjQiBlXrW8a0GtinbinwkhMhGlmgPewktVH3IOkGEkECxL5oVgc9TZ
XDiOB5gJQvDc2Rwlw9f6vWNK/5yc0fOaocG4ck+n1AY40WfBW5TrXawjmuStrDA/jGNOEmybKgiE
XAWC3JhbCBAL/7EhHUTHltBOLEb1CVchaBcBMFubmH1CON3eepY82Y7O3LgexZ/RH/CgdOpOA5mn
k0ZH4iIdjDTqoNpW4ItwJF2lCjAU4GHclbZy4RHY+d04uLsA4XRE3m5eZb0P8c8J7O3dA7XUkZCC
rwOXygFB5KbcdhnZP1U3fv+oh6qiocUrhute4oSfvmMSMBdQmi7oXu07ha7XyttxL+noLrOjxooX
M8VTAHQSEJzLmZuDVndBJ5lg6bgGDe6Hq3adDD30pnDMxdHjIjDv6gf0YdDPNYGZzJ+IZ/U7rbRr
X0NJrWxbFQBesbYMO8/9aF1u1yFnchG7JaDV9TIg7LPr6M/Ep3yoSj7VsUFdf0WVRQiNBM3wuU+o
RGmyPWTOerEU4afjRpTf09GtVvcmnGZf1r1ILvymSKFmrorUSvDK6aWDaclCgTrt0qNuopOsaVZn
E7dLpx9crcNoGRaQvpD+uvBiy7kzhJxyrUwraUQDmrKIyEk1zsMeitUi57P6EFP/G+/c34C96btG
g5KXvZeqhBD74I6ztChZw7iemVWlq/FBF76lq2f6/2MA5JaSDbGJFS0ZAYXvHq0U+TaNjky+ggFj
9mHPUVPpm1RQdt0TV03v46v5erhatM15hMB0KE5FsJlpRpZC5AhbKWrF9QTat1FjGOuILughC7Xx
3aERUBLAdlXLngiRapZZNu1AHOHlNP+W7tPYp20xzWmlESdRHw/F/1GHe54I0XtAXEOfHNFOtGQX
k2ewLUUC/v8DUUpW7JZ9qNKM5KOzTvOhodgQuqpvByxhTzG/r4AcF3Ot7F28tmRdYzabTn3TjFfV
NwdvGZfU9YHgAUJGvTOU3YIVklK7fWriEhb7kl/Njk03UFiCxiSX0FyQjjvNK7lKOMpO8roOSMjK
BFB3F9NCp3FpqB44vMtt/HYzkThB4fE9BFjkaBr6gE6ZopKbIvRWJq5Q2tNEEGcMwES1fkWK8jRE
srg3VLZ9k/GV+f6YFJePhRCydcOGGITaGb/e9c9HYOJCum6FXVVFFM5OYJio/i54yxu2bFkxds59
8c5GdjA8GHINf9u6kup5F6LHRfHYrpyK7cTzAGRejnuhsE4eCt0hXAz193ZTL9mg0fGRgvP1006K
nVIguVoIGMhQKFVeG2GHw6dG/RHAIlmwg2IOuC2RjHJcVWBkhXk5N3Xn5JSCMLF7miyiU7RA6/W6
7YhQrfG8uS8XeZDyKt2gV9r27I1bM74xzxnmQ6b6Y7XVefbh7viluFwfGsHcQZUgOzFxMKcNNat7
A1q9YIo6pxwdu42UO5BPUzEIa4GhrIIk+kizKQHeKYvr6vOjQ0jLfqV4RZPDzn1P1klgGLUmHFn6
cjkuS3Eza2seSWRtumG6XnSw77lcBjrCT0Y+21mUfR/2zo8HskFoWFASf4//yNSpigjAs+ADyiAi
z3Nbnk6PcEzpVve47glMUqnrIvjH5hr2dzDlOTCYlbjZB/l+OULNnFLIoj/2Wtw2aI5wQ0ua/bJ/
v3HOVcWs0XXAu3A2yBUsfP/Fh/eM8J/nMn6p/XZqgOuUdS5b/3g8fXn0LzLQuTCNqDYDcKFjuwPB
m3n1HGN5OeNISCBwwlsXU/LtvaPmgneIYRXZvXQ3z9NSsCR3VCQP+Yd4GCKRhlhToqvN0cpI3Hy6
2aiwNITkmlvzmumLo1ORj7Vz5fxTBgUNbhdNKupJhYi42rGCo25l1UPCkEejD5Oz7ZCMp2xJlbZz
cuRS8bJ1uhfC8OnOKTwuVDyQeyRte3Uk5g/oRMpbZg+CWnxj10ODpkq/K92/3N2cwfRZHRxXb9JU
dxnftBQv3lt4bjD2OMOUQdtwdP3astwwN51DBKihuM6lsd1iik65OAsfCVL59WXsJgaRObJCMjSF
XzBc40GEVqkNu5WytPtY+eTcN0M9mi5s8w/eByB3xmkxugiKg1ComTwO6d8RhjycnC0S7IE+DPu1
6lbE8OBuX3Efy1tXhcQ/cdDPYSjso9T1seIFxNAjyJAHzesQwd2+u30e48mqJLKX4q/mmgfqyMdZ
lL55L9zUyFi0ZAe/JFkCZjjZ+BegK7+8fm9tNNQENQJw3ij3vPMDBMfZZhtXmgxrw2FFU20NmwbB
4EYLKyTdMTwx1KEbjwkM/naLP2ZKzKKAh8jCRWtWny4SI/X7HpQwHeBSgucKP+5v83WK0fkuUo0i
0rWzJeQooUMA2pIqGgVV/NyykVomuceYEFRqLDYEeupgtt7hbRhve2qp8CbeR7310OZEEQcUBVHj
NFMElA5abz/uumVYVqOSm84GEKh9s8+Ei0QbLPiBGwHlrdbEu8h+F0ZSoHL3uCjIrcG6JfveBck/
w5XhIi3Ore0OXRldBp8NkeCnuM9Aep/J1fdrS2NXhH2LPbzRMxUXgXgyAUUl7Xn1zabehrovd867
MHmaN0/JR+ejKLQRSPM9+D/IK8nbmxvlhIav7Pas7ccB9SNSTSQCnNhCcaa1SI5GOKthXVshH4un
3HYIQGS0rW5HjBO9iTrreV7X63uQAX4Rpdqv1++bxJRD/h6iFihQLrP0P2CS+OujkM6Wap3MCJCv
N+NqQO5JkJJZwYQ5fd79I8g9Fq5eLl0DqGOd3juBAfPjk4hkcPMht1IAciCXxdISUGhNtOIZYDLY
iQ9qdJMjBL+OAPAu0Yq9410NFPCkvWr5SWRlqq0opVVmVLAFPP/mt6i7jmWHTfxGCxHr3Gk8B72H
SFjV6AwZBk4+r+KYtlIUH6K/cWfMb9kZqjO/r6lJPhCPfNwGbIciTYCLxydvRCFhg70naYtkkzV0
RyLbwJh6izeHLL1JzGMUK499P+592aPTZAsWU3ESGuAFqS/KRO67EYvQlbol4YJK60BLxVPR43j/
JJpJLTsi3njerT07bhhm3QYdzR8nPlcKvBnQXMCnkfxrqrtc/nPYxXuyzQakD9FmZcu/2ssOvhr7
iiKpOqcM3HXVuIerc4kOFCUatuCtzU9xH2NRBFlaLUl0/J44mQCpIV8tNjtCgrOVYby2ooIV7rAV
IwPBpA9AMhQL/UQWq/dSh4VK6zz4oLS2dM35dkZOTnB5CK5Yz6R5dPvCRyIys6B1Lklz3Kb4T0Jj
Jpxz4qY4xanAP9wJDSHlG8ThmWgTkqncbhGYsVuHoaNqdCvIBbvd8ud0+X4d2dsJXWepRJAH4EmI
WwN+zerR2WaPtXMbkxzJl9GFJ/gTZwm6EIWG3TRAiR/h3LryKdSmkpucsG4p9q4sQzcAqn575R5r
5bkFCWemWoe7hqpY9i/JHpVwOw8jBtridngPNtokLi9m3lLnLUcO/6BPY14oUovhvcGi6jQ8aIuP
LtxA5hWyPQswW5wLphJebT9FfD3+y7LPXZmaTmsHg3n83fbfcPhmdyUpaqtgUzuBBdGa1Zsvi6eA
uHLwJmZJ0ME30n0yECXKKOgzEJghAjpWCY8WC4MAvPpJSeZhAzc4aDo/3JFTnTE1kTZaitN5vAFN
74l9NZfmSuJ3D2d49tEycG4Kcqk3xbB6pdL3zuqhjTfV/oOKtYS0o40mSGPAySe3WkvkEsTEzTO/
PseEp2LPJmkWLyR21PrWXB/gI3LRd804nKUp9eYirO+HQvSVTWBX5+rpYf0jWzpZwbP6O9Cd4PcY
4JPRrn6kfTxksG+dKDD9CRCqjMbb9c2oOmq6tDC02aFAELO2SJ0uOR9tV7yzVLOS6AQGD45z92X/
epVBANoraGC5ZZhejKIsaniuspZL2i+nggnFQBzp9p8150XbU1gR+gBH+4iDPF6ebX51+1nhVLN3
6r+jvfyzoFo+w6gXcmmR4HlfYwKfC/Ts+pyZ6SsAQknvM7Q8BXCHqPnumpIW9j27t7GkE6WnYnYc
Tef6dfAgPPAaZQisfj9DdLJvyHU34zTKNkZszQfXe4s1+fkczzCK0KN+NRymCE1GfoHWPMxy23CP
jhS4gGAWVxrH5Bul2wASCMX2R1XuVRprN/OxNSM3eZixYSJ8n9EUCNIhYMO87hPjQQ7WUkG/x3z5
D/JhJGtzVrhm+DivEjriBODX9TUt01BC+fFhx5fWrDosZt8S9LhkOnWyZ3fmE8NpCBumb3rLdS9X
Drwws6HNSSQMoha3tRcy08daLLU8FJxuc5OG5QoXQ9rJloFRzVAJytuLFKmDussRY1ii3h3CL9kg
Mse8T+yP30j4081QRJxVFnlNk9ywdKzHe9mcHl6Z5Zmv6yCDtRuQ21BxIeEZki2qDS/IsZiEA9nI
fkZeioDsInpXxT2kGWOtHA2MJnrgRnPsCmfRhixXjRDua+rPLCGiE2oftk0m8PM9uei6BE0WrJ1W
UkX/gqVQfwT/GXRhijIVwaUNFnkvevjpCDFyhOrhE1GU7B7y3nVXQAooafj4c5STvuDebLFenH7a
+M7ZPg9WTMBrWbPPPn4uAgbbpJzDpIbwJwFInNZ9qYSD1zLXgVOEkL5ruV6Z3IJk/z8Jo8oufMFg
fwsZJFYrcPpVmamocEh7lH7WRsx98yG0GEXXopddYMJLZFeJ4LPvKy7qFdv6rQ0pfuGJXI3+t+Pf
TgbOhOkuOerf2WLRxBJw9fWBxxj63l+39BaWFouGO1gcEt0XQhP4ZQ8cSJ7RwX1uBSw6y3nJ/mmR
gPW9SePPj0ECMGlodZMEp52YvR4QFXhTbG3ppAgaFuqjRZpi8yVtCwrgZQcYGt9rct17GhbCLmcZ
E/U7Pskmonj+b1eP6K+COZ5+Fe4P2A62ld4njpZe2jwQFuVfWJYBXsMdKbA/mYP4IORYRpC0Cx4L
MlBsRgIeX8z03M4PcmTuMvPwTS4hibtav3oXr/06wInCtHoAmtT0MPeMBLOFk0yGc75+mPxRIIpw
EuDaVxYjK5eZ85rWVlx9wLGcxokuwMjqd1Vaz0y46N9RhvvWhMOz9SLoQ9nH2k8iW3q+NBI92VsH
wyZcLyrDz5jXCOFpP5jgFri6YTw6TLmtbHsXIw1eNlBYW9MURO2dOZYSy9ZHE3g5mc2x3AMdhveT
DlGdeJ9Rh+eaohJDQFHlahdnsPLrI+bqrKYN+vxtRWGucqhfrR7DdmIjq4virIei+jAOj6Fntplz
Zgz/2m4PYvGQjdfSRxD6itXPcr5Ts/oGNwe3GNtZ4hfdpt1CFLAoN7RVoyZmy/hOR0m/Y1Aol1GS
TfwizetVDi/TEiotUFzr0FL2J2uTztKDeD9PhmRPX2nfczKmTQ6q+wE4p8SA7WXLeSnDomckMqZL
8x5JzSRhjRewXUPTH5mH3U6vAsDfLMSiD+OEhjefMyjtM4HRLafaA5q1Fg2v6TO3PA8Bc8p3WKKK
vawsFV2G/Rb7gffFugQTy2hHHZcE2YLmXIr65G5ZWlo6C8wTnGoiW24v8WcspQlqTdMoVve+03hj
dAs7ZohfEFVMtfwUGC02HSPurQB27NAUAp6OtOgTLsN1GatEO1sf4UAmw2IGG7FVamN1Yjgn78vu
Was/kQn8qFoQ97c9i6femeuY4O8puWFE3ftP23XqyIqtc4DSXjW1SaZbvqEuMMWT9+MfPHAAdz+F
cqX5qq1QYxV/2bb0ti0F4Rt/sDjvfpVPgFe/ka/qyo8f6XtEImqBhThLqXM/RXq4V5oRRyWntCNg
BBEy84wfvxcVIEeaiXyFtO9/16TQ9wvgoxcvlZ8ZILtQQ064thd1507MrvFKvt7NWj4IVmER5LRl
zA8B7iFpN0tcJqiZZmk0euqCIZ934KECh3qXLXxzD+8pS3bVtAJw8livWEJKJVgBwLLvQ45X1R1+
/5vJgR13EZhwl29+OR+c7CI/J1qT6leloNixD81WEj/nFaXRgHNTOUE08YHqR+lXHR/Huik134Ll
+s9fikeh9YyZXcSlzh5tjjAJnpYT+sUz25n9S1M0lZF67PCviopOAJqbEhqKOqAbYeVifEHcY21T
/D2NyJohs1MfDWTPpoV0cP3VRiK/iXYv+P2aHSplIJ3KXV3ZXeQXxU/snB/bGh5rA/fnslY62OhM
1DEXnKxk6P2zHtyGKmDyO/5oAQTFWscqhHiwcgGtc5fkpXcObI2KabD5bJ9k84nRNp6QB6EgH4pB
Pr7K9wS6BcMH9Z8HHQZmxfn2ymKw1bA2XGOHHMGm6ZjSOQLS4+7+mKQSUI+4X9CzO30h9YvdS2x1
aUSFa++bubNBGkknjBlGzQM6GWN1oXByRqsQ8whqr0NhjVgbW9VdoaQJ0YnAccMl/e69NpbEyCc0
njED9kip6WISwnx/ry5aWUZZg8Q+2pHH6vFhvq2AcMpU1VtXhXMyBUY25Gc84j+MPKaviJtH3hd/
9LbruudZGFWbm0jjAHKFu/i+OKLEbwPqYJRbmUch6ZxMfUNQSIXc1uqdH9GtYWWpiUyJOlabzVJ7
87Mh/eQlFhHdz94WgAqxcoBztsr/4WjUchrc8j3pGnB9YMdWiXQsBNA3eF9wF32ZGX3zPdG7XtjT
T0+5fPfykMkSpzk6bRo2oEoBxyn/LYE+djQ88l5xGxNC8kAG58MU6p70TT4Tjiz7AGZY/xSB5fvi
+SpXBwWb0y0ggvL8Wwyl7TFRFdFPJYVSOeSxcN+mSUJsMrpPJRVHn2gqZvkJDJyfZhA/bnaHibop
JbVKfVTimiS+GnDHtmAwZ2DYZcq306ZdqLMmbHMaYWSrWPwGbNJ1l1fkDg7CQajm3YSVuSVMIQNq
DZ8WZ6Qp9RgEprg3sC2fpnP3bqp88WAT+gXOI+0PW7fuNlCBpQKILrUfnBdRB69HlwaQYHbBN0mW
GPk7XOnvroZhw6Bs6UQ50+mHfiJGQ1l8gO2VDIcjH1cXQLEoo2l5CyY2iBxwlByZTKWWjKK6cbnL
Yu4KtjvuM+J3BJOLpCvze5aU58WTdpFsmb9xGYcpxoHEFZkUnRwkI0JRRwX7i0lQ0iut5CFOqlrZ
xoKzV5pB2Tn6Fxem/pEgZYHEoXdlvRAMyqrKPFDjR+eVT+PCFmqoxiEg6IZp/okHQ9IU8lUFDph4
n8wwLEEG9YSi8B35hpL4r2pQOM0kdD2qUblQZmQLn3yvmw6x4IBzZ1C4Dc3hP/JCjWjyWBJPbqt7
P3suUdReCAWeIXEGz7KF0MfzRpn6xyyaSUbwUI+wgHEF6zLMqd+FOoIgtR8TgwpiN4h3AQYGxVjL
emCMKyzqce5NH9Gl74buQOIwkXP+ktBdJISCRkW8ob28ygV0lgklNjV/dHbqgxp/uIZBTtuWqAiP
KWWjn/yjSvXu17xWbdd430kMOzFOH7YUcGrXdX2BIGM3H6dJWitBM9AVrEH5b91BvcYLoP+QzQ/c
xiZ4qdV6LlW4tm8NIDmQbvdIUof3Pf4+Djg9Cwt3wIMETUsWeZbjNeofgPUh4V9RgoFk9pfP32hO
4ZuBbGJ38rPvUyVVheAQF4m6R7mrQn3QR9ewGRKewN4WgS7Hpt7RRrZvjPEBdm871gf2PiuSPi0W
eSNH5sHObqDiqJ+jTlWT0/HgAj4ESZZuMyebVWaPVWGDO6M1NuUHIDNuAXYKqkXkLDvbrlsfsTc0
qOICNwWQKqveT94UUmFRSf3BXryf2iH4hiX2iVUWPnLij/G8b62w4zAIx6a0BwPNkLP39VkHKXCl
ckSVZOcNDFeEJtp5xjBJvE7dBLlOC9XsafYeW3SbkqbN1RngRkQb+d7IsQDs1+BVrd16ZVAr7ztw
HpUlZsxwABmunDp/ghJXDvaH61yh8frcZsWFetrTVQVmHo+Vs3g1sUKxc4h8JCheT9n9TgGQnn1t
O585sVceEUqPQsCMyJXHY4YmygTkf6U88nDTwaEZ1bzZKmqMIKg4lzVt+tLtnvbho5qnyLjfcqyi
p/uRFIDwGSrHf8segv412HXoTYLZRHdYVTYIXrdbjSB5nPiEY0OIE2QH2oV/lyv4zVIY8+ctZzzd
hgrt1GgC5Q4FYcHppv8vY6PALihOtK2jd5Ku5MjrV81eFlD+u1XRhthiQDJyzCdBM1NFzz9yWLrd
3UjLwoRj7xiUOQsG8hukqt8dRfbLSd3Jbsc8HSHcmGupFFgJzbXQp/JV9QDbGMlufhGefgpI5V+U
eIpshL+NSOvlDwaixHugHT3e7uHp+kRubrq1dkchYPUPd1oGwcvXmT51q+DOU7JkcGQ9lqa80mzC
3l4+k+Owg/HoG5il+rolnwAro9eM4k5DuFu6dyCGAC8yPIrnA1R9R8VBD4fP64kTsahhiJOyLw22
ynedCHZG/vAGb0qxx3KYOWamNj9zIPjgTOqiIK1fcjXe0AQm+p3+sMIZMgE6+1PDLSfwb8Slg0hh
IC6JbkmFUYKmwqR+KPhrBmDU4wCnNZ9mu9FUIgQOEAAUZhMCwqN/HORE+bHkPxBq9aXFhxxiRoZf
0e1lQTTXfK2/PpttB7RFyF4jw6WMLmVBiyYT4Xya4oePu08zRDICyHbuMhmaLLzvSARQsikdsNT2
M2KEOX6n052dWQL6Yo/VUKVXasXcwikThb6wJuK+Oa4j50RMTVjGnWcQOYyBn+OpPDwdzPZ2dFzi
6XoBH/vXuPEXlO+pQeLBeVYIUrWglSSKKwP8Y45OJHvF+yQVTOe4RINPrOJX6F6Iro8/Eph00IgR
1NkRDHWxXMKg4uEoC++sbLZ/Zq58/oQYBqunxnSQncQNLtT6PDkMWuF+/bGQGgXDeY0BiaGFFyQf
u4nsWTWCGR+gjEe3owIbKHVz4pG23E/LVWor+RKOPV4M3db2QSQ2QKAUC6g7YOLOnQFR/B0WO8I8
/lzbF3LCxDsib6dJ9ukbEPtPWYm4aAauemhHrM4IXG1ziAnY2GrH46zRFIag/nMijOcuKkP+EqgP
XXavZoFV5i9vv2wddUV7l10LrHueRH9wMnYu8Ruhg+82lJRM3QF4C23WqkgwUA0tQ5TX2fXclYxI
7XyaviLth/bT0AKtk+lLQ6+y6NIkimTscLMmusUpXFIm8tfAbR/SzIVpPeA7ql0MPFro98cMSQiD
UvANyrrQoHAlv/qfJcURI33HQVZGM3sH0fvOaXvZn21bbdq9EGog0IpIAEgguqu88e5lZvfG8//6
QGhYNhD8UxkGkju3Zi2+JpT01LyUc4CzfrPbcw9V9X6VNz0c6T65bLizqCVLb+F8E9wK0rTsZFPc
baygnkiTWooErFcVZGlV8eoKqR283HxfTXRqocuRjoYUesPu2xav/3jEgaTUqqn2nRKLZIJGMdqx
UNAnT4W/RCcfB6V+KGC//UZB/4GMjjgts3odFlPy+WB9Tsx+fbiotzsk/Xpgi9zds3cFdF6VzAlz
K9beJX8ylWx8c+D2c3XzYx/N+d/N3qpDU87jJxOrmsOZt7kB70AlJCAP1tIfWsfrI+/zU3h+u6il
kfmBTKoa7HbDv9xzRKcR3t+b0grcmB3A95mbQ7OjJImRnGTuzjHns1Uf4yu6+jPVSC1tiiXWm55X
7qCQytuwdUzOeJpaRoF/1FS05110UO7Ph9+Nmmn4bYZ/IDgbtPcRPtudemyWIph9/1dxG/Sr+dF6
IKTlXHZPV/cCzlEdUJQPDBgMivKDFUdeW+PTBc1NHx/zv1auxTYS4n0DnDIx7UyqbTgIMz2eI+55
mhacv+cC1VsajM5BMdCc/0vQ0KEo6FOU53+E8Byxc7n0paNBO0WdSzQtgfOJ+NH8O21yN3TLF6OH
iY9qSiBvvwLDwgumnH1yg3Xatv9NjIJe3d0O1p4bB4Qfv9tuuT+IWQrVqlbW8mJLfF48ykyFhQuv
/sk4kuPOCf4NqyJc1iQoTgcdJ40Y3XYPwJI7tlOB/iUEEiw8qbNO3Wuk3XT1eyJmSCQ5SWIbG4G0
uvYvS8R9Vavzl7iTrYi2FYOd/y1PuE1ULcJOtc3Ln/cXkqxW4ixQLI/XVT9XuKrzUgpIePQJ6sJw
CynwBv1sXil2VCGZMNPsTYGhpQNHU0JXdrR46tMnvb3XoZi8VexX4Sb+/cX8mX8Rfn5MAJS2IVRo
lK7ZfkSaXQyuzzrKAt1zNfPj1EtEa/9WkghAWuF/MBlVDmxX3rZJsoM8IXCwBKDQfHfiaZFrcPkN
ZIXzGT8vAZv3/+jt0fF4fAYy/p9SSl9DxTsUG+tGw/VCYtYPuPdEP7kkM7yqOejT0bPrMarA8V5c
hXGgT9pQTgLEMJqnG6hNCRBr6OD+mEJ781WXsnQt2Y79aPNSdM3lCMTNeXaMU4Cd1vyiqmPxICjd
OefVjcbwUgI96BajvVgDuTWXwn7U4EZATz2kLuM8/Yni8mIPOMpA/ziU9omuGjPOYfrKgM8fX8oI
h8Dqs185rTVhsTAMrVHI4uHB6ba5FFuU++PUd8tOA0hsYROjDpyxPQcXuemzqDddLiVCbRVjvXo9
P54FuL7+IEOcKAwny2cEFaZM9l54Za56SZfbntYkBGNnSjXcMUausPuXE5cI4cb8kzVDcv6NyDTG
Gc8cJYzIvdYF7T6gi9C8cDUOjOx5xn9Rg+dMryNSWHjlkkVn+SsT7Ymn9X2fs5PLeybgiGas3VL5
3Bq4uPUzDnDHGzse5vJyvE3LdFmC+DoVV0lEJtN+M73LKkVeqy3cEcHo7yH4wYopcJHc6kWcIqaD
xN+6lTCBjejHG7BCZp3x4PwH8xCc+5sMbMAtNtkEYXZ5f9+EcU8NqLk3SJhTc4/WR24PyxRaq7HS
A0gPgmQz5LNK13DalaNaO4ljR8zofg9+aGV8LmJ1EGUXdXrq8pDgH1V9lgN3WaRsIEze9DleYa4z
ukHmXRbloFR7duHVCTLTp0jq52GTNd9a31bxUBCKc9HeHVRnhpauyblK6Nt5A/oZSE9Pba/C88HD
WryZRqisVO69PnEKRGiDDnXH5p1QhhZtwE+Q3R1Ad7UfH4cukNIyyrN04M18+TE65INaCFL/AepN
Xt/LKm+PYlm3qK3sUck/+PYps5+Jp0zWHYOKFHI6/7RW8EsSKmSP0vRAacH/F5/a6GMJCZbIHdri
vL4Yl1CRXAL7G9Q+Vb2oQ+2lOf36/6rxyectF3okz0ytx6Eqk/3GQlxufASH9OjMwYevJmjtSJaZ
8Ifg1c2uPtXtqbTYcb+V65phCCfJM7vNSQXA3OukHLQWLcLIVRMTIRBJpxB5NSKQEuI0cz9AcjHc
zIz2oOieyrbsQBpBpuFmuusxHO1Q5PHOWw4tNGe511whH9t8eFNhkSW/rabC1HYA4O6436WhQnun
x6GBf94UdqWWibnKLu+J/k5zWLsFq/c2Oc3jVodD9JIs6vaOHVuvvTHpPHyA31fP5DE3fRK1rOoQ
/CdyOFBs2GfnEro4jhs8im1sxbUUWYO1l/SK8ZRpA7XaRIhx+irUp6BbCV2xwfJDRwv9TNIuOn/6
YMJtppHQtyFtDB+DQQ4WPNCjUUg/doBLSCxiASXu546Hjl8hTcI9dWLc96rP+xAgIOCF+o4yYIpD
5IT27yFE57IAaxKf3n9oa6Fa33nt2ayGeC1+3N/xvMbDEmEoseI2vgWZzGLeI8jEsAgfSrh4LOYS
c9HzcFK/oV2XyYUaeV/zxt21ptshae1W+j26B8PQI1qpAn2R+Qalw1nljpD57orkXZy1AXzztcaS
+jZ0IX9U4+6nv+Io3IdqHiSSPRBlH0TjthIoe7RWJ5RZGK+011DNmJfGfpKFzOogDDKxkGTlmwmg
GujdPMK3oDkKpJIz/f49XXwf53nCJNZ+1uf0gWTckrrPGQctnOwEcAygpoGCe1TgIsKADW15coPd
SWmCCM2ySvrgN3ErDvxBZtSvTH78VzCbGlOfoIqiNNddxr23jbiKQ7uENxQhEq2Xxq9mGAX3Xi/Y
q2cuE/z/TQh2KDFfohw/RH/wh7bXdAlr2U2w73KcLAN9Q4/3zvr3ugtDvR/WPVKSsSCKEn52Ag3q
POR1obkYBnlSuTRxeWVelMzyW6ZLAzyXK0TD3qJg9fwJKQ5ALTiZOd+OPuZFVfxijIUnfBpuyGzE
F4cdyZxF2X0E2bNsDJ5uUftOsdfDUBOPzpToRvl3ba649UfmGgEGaI300LW1gIdTZcxp/Iammva4
T69+JIiHnkTDL+YLRjrja7s0iTSIlaIJMndWjokscuzyVWY1SN9slU5RumOiwrth7/G/ClglAEVi
wGP58dr3WiMYDhpebPJOzIDp3iP1fufR/otj5tpONyXqbz1cDy5LbAOCy7TBK7rwvpBoQLl24b3r
C+3hNRF0TVn1AToNQ8M3TYGsKhfJO0kyuMbsuiZcyGSHKILwxPSRnEBkFg1wD8SuFghphuKC4NY2
BCGfTsqRSeIVp/JlC4FugMyyPGErveNsfUgz8fuEG9fKcBOcIPrpJwd/LU1UCJUvXGtliJCD+rUS
Jpixve8omc8Jbwn63QjaXsX8R0tdhpB9GCgy0NwDxawawciBSp0gv4u5pcovUcj6EDMmGaHd4MMJ
dpvVEbiRPHOhQliaKMLn3Z5DdutbX1ip+XcyRUuf8j6V0ovGUiVJe+H8deDD6qfQe10AKfr9lvsy
zzWt7c9X4oVWOmt3UdxxqUlLP/oj3S71Zd8Al7xvR9d7+4GODB9TrCauXl+6cxwkPjeyeinC29+1
uNyWjCARCuCXEV5VaE87sJxQEpoR/CWmFEVRsg/QMdujsVGGABsNrpcHHt93KOiKPOe9LSmFj0qo
5PXdONtTXTHv1/2lJsm0xuetxal757XF8QPewEq2oECBBkXBTDJGxd6MvKaQjkpaQAySWjDgfHQG
Bd9WKMWXAziPgOnaQB1HtOl6ku7VNywfk5pBAtQTLsh1cN73iDgxAKivdBadxZwQlH1NMphfKjgi
kL81JljlPD52HrRuE8GWIor1C/NGT98WXqRhwp/t8GyIqhzHChz5wIMrI2Lw5Zd/CdGtQO6f1ZIn
zyN5wiNSmASlfkABQmMmerbKz1V90TebJSTVWTlu4Wxvhrd6HcWRRQiahOOEWc6ND+OtKbPnUmB3
ZzBJFnQ2ZAXOT7aG3p8HrQC71oGkZeejqrt7QQyzY9e5vnCUwTBXkPwKMEeO8wHx1GJJrsuFYWBA
avASoVoo1GTLZGttvllBW/Uh4Py4m06zFZsBRrEONXz+WRlYt0MXb+UE34CunRfvvjTa/Y5bznzO
FTkOLmxNrILVm8BNCKi45ZR+mlhHbhBKlYdX102MAe3XoHz282S01yQs250o6UmJYAYeiNkum3hi
TbVsSNnXBPHJF4/IoqlaEHE/oAybYt3XZ/xqNVLmeWlMCQNcjip6tcYn3stxTRunQzOTalGk8xam
jU4rCAV5oncA2aCuSF3/QpiEvGbDJYTNnh23q8qGqt4zBnNTxikGQsFXYRjbx880j1KcN6Q2ajP6
A5h3/E4O/T6Wi8NXq1pk0sipOXLV/U7/tOoL2Fzk1IjUjgkSDEafkjKrkt5ectj/nsB8uDNRLJIw
pbpWn3ESK+aCeWBdLu6BNLQMIx7gfMo4kb1F6CZCI1ZMsXAoMaXvIyY6+fh5WwjI+Kdnv4QlSSe4
2hmqiYt0cJ1JwtoGGGEyuKBauKTH2AUyArzOXkCnwoCshbUriyXj/2FBkhUDdvvmt+nM/oLhg3wx
jc9Z6rfeWpj8qMl4kQqflTbHU+v3Rl5dsti2wkA8dTrm+XLsD1rH2eeXCs9wOhyKtcmLhYDfrHx3
0+Yvy0ZqbkXhCPXb07cNg2nxA/ixRRGe5N7fewuIdrZUUnp1Z+KY5VLZwEIGr+Yz8cCpqNXJYfGQ
fwmJYokiINjMLjQ0Q/ZSLbg8npphD6pbFG7gyWG8MFhYqQHnmAEKrdKnOvP5dUE7mEKeRLijCYme
4AO4qUEQkAW+/5P5P7J2Rjkyz+lfeKM+G7/lKPTee7fYIp3hhdJR4/3kMV8ILZ5s25CNNcJa2ucX
T3dPEE/rU/hzr40Lz5X6FRSasijXxn5e+iuDxFtvzSvB9GjbhF4iCRaFNAUNxzHIxiBYv8dHC+yR
++uD/HF8kqg/ym4LtDJCprPVcd+94jcdwplu/y0SfYh3jFmXwtSb7gfPM280J9cDAtWV5JaLQSi0
h0lx58mWR3tfs83wiCdpWHbc4x0b1t96o7+wmj0/rR75vjYawIOZiEUamdBlHtmdbzuE4IYhcIIY
k8yBDJmGiMEEXQUV2rF5sN1YE8SUrwK8vR19YeaYRTlZQTLb5XIEyCD4upVX3GVdDTcCFYloomc6
/e+X7JQpkWqcX1grM35vi8GnCORuK4LmZbu2/5/NzYsuaFiAk4H0Gqp+BaLfyjReS7YgqrzDPJ7m
VtrtZa15F/+TTptVnxcD/sPU6j8PYadcNV9f9gxoXbRK2yFX0TCLuD8/SNjJaeN5aG81qEqOMfDC
//skXEnZPFfeeTnTOrzOijRQLmZ6nJGPeC/ia5alsriXeL42ZODA41QP1ESf15sNAc8/+o4Xe5t2
Mnnojb3HFALGN2fJGVY0DGzVhO5NM2N6A8LUp15BpRs2f+RKBG3Bk7xE3LlYCGFf12FWlK+TdvJY
aNpTq2pesu1EgRNdfd38OctUlveM1XLMIPFGM5m84+c5f57gMN+/1eFUKC6ErcHZgBawTkllgzWv
eG/TyXyHlI5WoZSfCEktNM2Axxivvx+MwBAyblxjiQk7fWgFox2VsoX6aM8VauUlPPDONgO2Mqwo
jxUvZIxRadnqrL4qOYMMc6ZrYvg1AlvZ1LgKKenWoT4IMZWcpQ8CcOTQsn8vE4i1/MDRnrLElpKu
JqtzPAussf12siugAGtg/qtq6q2iN1MyOGKqgzrRip8nje54p6uCCOWt5H1IpB5sgqcK8tvpb8ow
BExBeaoP6izI0Ghf7sn33BanGcguWJYCFSk4Xea6+QTGhszkSr3NQ9jAmmaVXzlFyFovLSn2IOET
ywG0BEH2s00GyYgd0SeTyVr/ywPcjfXL2oGL0nb6t4aWHbm8bRHTKl2OO+PybAD0KO5L90BJZn7/
nwiyX34tTRBlXoi02JZDPbco55AcmmZU2na+0ir9CYou8e1tHZOTDCfosGpE7Iz3/tG+Cb7pjM9q
K6aQfBa2tGucqFiIoI6W8DKwQsIYjgCO32JlA22aYf4jlYFq+98WWLlqxttCnZpIG6znbTuEBotM
F721nmnyZ8S/8olElVXzDvPfP8c6Pq14WC4P/WywKqZhIq9GMsgnwtFYRYA5dTNyLRkH1CK3NTb+
u1mc/Chonq4/cSWAb1NjSO9bAmv9LZpwnjDTS+d5FwmR+2v+fyQGWA++bSBuX+rSwouMy1Zba7sw
ZPxhByc6Af503eQwersM2uIdQ7Zuvr/XSlBbWelhv8+g4nlXesNOf556EnEPSjr2rv5HQlJCoj17
SCsTrtWBgWnpzE1pHpwDqrSTallU3pnVk3gNtEaKpws7CGHgv35ovbvnoqk9fOOC0rKX2KvvtTDK
6KHL/SBaKbmDBNztXcMKwd8kGA5mLmG244YxlqzKuDLjPLNAXlKciokao2QUm9Ftsfaeep0GniYP
AIEhMwc3d/vYYb9jMk3JRm0AIpaNu/qBATTAo41zdEmuLpqx9Tcbs+OB6IhWXJn4fKcP8WffqL0W
xrNbzme75m/2BUFZSbJZxMgkWwufK5rIkteHft3047V+pfmeIW8jEwM/x/lrgcsnGD1UKTQULoXt
UGtU65u/Kp7f7zwHXuHzxq/g5wShZNMwclvLOPB0if2VRmx1Og5eewmrJ/5aQ0NUmzgt91dLjvzN
3uU2a0vUZORcfhx5nMa8XyXFKnGZERxb+/rGjfhPk+l0xNsJ7oxX6GzkWt3RQom3OVdaALJ4fFIK
44KQ2tuUJcILb+R+CgjxTRfxF/OkA0UGejaUgxvMpes71y/4M62hlGi162/5831LXGkpJN0+7//z
uYyJ9T11D571jXgZjCmjBmBhFy45Y6wHJUyX8KO5h7NtdbuSHOb44tYn6Ml2kF1hzSBvJ5RcjT3B
WcbJD2/+tzsPvaL3W0gJRZ4paSb4I5Oil+32peGjSjuik8SgzyAod2nUtxVuZK0Y+az1QO1SyxcG
V3/0vw+EarklVuP6Rf2LQ2CUNW1f5nge+RzldlHZrcl5HIlWkdr1F+dfL/PYn5Fl6YP805oQi2H9
AoI3XvcMp4i9KflKF18dSMfIgZnoYyXQjyLjjgh9sbJZBmD4b/2cG3e5zHmWMHGeHyQjwTZSaFLN
zFnYUi6GMpLAzoDAVXwwH7TlLm4eZrp9kNEnegslL7iCFs3JJedEhBq22pVOM9EpJh58cC+CdFbI
033WgI0BFUGC1NdvJaXnp+2Qzj6dCZSFoPwv+9IVO766XjpnBScZN3qDwqjLVs41Ct5aNPBmQa1n
tEmMpzHBZyMo2/w/0G1AWY/4d8GYxFWb2u9YdQIFCdLfZeurtGefmJT1M0YjrVgqfg3vY/EFmKoH
QzC+naNINgP8hfinzsivqD71PJRnOd3ummckb09QKUFGeqlQObfPV6gnxeGILXrum4QHcxInMua1
e7uystQp3K4QgEWQB0COzGDaYWAnIPeL5rTGNgUXuKYuxkcFhxaFsT+wthxB5Mc4+Ks0aY8Cj2/6
+5kzeMiCmXWdJSCqzBO4k2elMQ8idVTLG+YeBJq6v1z/gnc2NS9l1Ior0HoKU4Ig7yQviCXS5g5Q
hHuqfnCk8pcl0LtdILMzR8I+1ithv7bPae3IMrMtGQfY9vJ9QrxW4TATkjVNpJFO2DnnHI8HhUL+
aUTXdmT1tFQ+r2yOgr/jQPx00+5KBLHwl+iZ78UB/gIuKZzUHiy9t8Bd/5gyT4Q6LXihj4iGFvoA
CVySvIoDdRMcGn3wmCdwbPM/Xhr+NXKbenUpe+5qQrTAem/m9r9rmn1k87+3Ttd8Pdf0LQBEiiMH
9xnrFlQMYiW/4wtmTkP5soLtegzAQVS4tUGBCdwHxaVwk18M4u7pjFxvTziWOsaP19Szi09wkVWV
Fb+WQKbT9xoCSC0M4KZJScFPEKaOnLO8XEYJyRoq97/y2/VXnmZtQja7EEqtLIq2OLbeEUqeedtW
WtAynBBzv1fKBxm8QVj4tXHU/cvJa27m9+HI59LDGhHbA1/nvjxnveJ2k23LNvD7udLLWUW/gM4D
QqTsKFrmq0ISF+SATCu+PzYh4s+R568cjf+SCwepfuCJvPBrR6Ar4LuqqH2QB1rKj9wW6bpWBvy2
aq7RFi+RP2/zC1p3k0KbRgaYWGdFPSwMfr8zNkK8B8zbwu2tJnaqmDYGQ1oOM/Fpw1jROKq1U1hQ
YD8mA2szrHhHauI6EikPrjxsyevMPJpPgjbj0u/CLpw5mAZ/bqbPj4c4wzCL99cIZNUDDXdVAs4L
45oltmZNjxZfyolodQAZCAD4kbsrsjdLt7htY+Sg1nF56ODHHs8vucnLhXQ0Vy6XHFusSKXhOVgD
0LG73/12YLz7MAluURoHAxSNLe2ee1dUaoAlE7wsDrERmHa0qmnGYTGqYwWBKJZXDoeme1BXX84K
FU8I90WqfJsxMCo5ylxU12gTjhzkaB2HPKAyvTNIvqj+NGr+dqMH//P+6IIK+mM9p56OXFDNk+in
pEDYuemS9qpsRw+v4dqDdpKPEJO440pmdoRTrH00sAAGaRuEZhcdUKic3ekQyg6I5DTQcrIHSWxv
V23FIl6VB3P09iPeRnthJUrM9qwnLpAj0vbKpgW+5e/5adrkRf4uYZmnH4VXaN9ztvtD9d6sBB3N
qCF2uhVpvzREhJ0YwenWt2S9VLo7c7FlvtrNG3q/a9oPDqpcJu2iVOSfa5EDSNhcUzHgNtof2+db
eiLkzVtwWXEmJF7fXdqmLNLn3aaT3eQeR0+IRfFCOSGv3LRATXwpDZ+YLLHqLDMxuxKD87KI00y7
ODtmNNZOb9n8wSxts7VrbFnVegv7Ygc5uvAL7dMcGOdyXDZrIVk5FTkbTXihk4tjJUHoxRHbF6uX
JCtadPkKAYYxOVGg38SaGR2XAJCKo4UQSYbDI3U0ZlHjs2LumnxX4Uo9WSnLQ3d4JM5go36HnMCc
yj7y3iJlvzgqXe1JhzFjk7xviyl8wYJ19LfpmBGygYJ8KsyLaS2oJXrlig+qSh8rYUcnqkLYKOod
m9n7iv67yjwfK0dpFy2NzKRKL5sxnufxHTGT4d/P7sqLcQxpjwydaQgOkHr+TxwXQf/s4QwTKC8k
+pGoZ++8KaQTiIgRFWSqfjXRHFMcIvbTjaJHMvDG5fpMeZ9G8obCljODA3e1OhemRJFfWWSzah8Q
n0fm7H0aGnIbhk98Nzs1VTNzT93VcSrqJ1m5DKoumi6pDg7YQDeI/hnkCMHrQQEOsxcLqQvqH7/d
b/fVf3R2oZg0scrxcQBlYJS+BUeNOX24138caIBkdQ4EYAcOaJNsXEW0SHKk+IfhqMT9xHS2ccSt
4d2umnSoHo2XbEvlQ69q/wTIoBEMpErK9Zt0j9yZ2qTchj75Jz4cJhnjx9zrlJwr45RWHv2eSTgT
8oGwUuAeqL2/lmC1J+RBopfOxCPOAY2EMdlKv/SE4xZ58WJo+vV/7rXfbsVMyBeMTWTPrwu/kJHr
RvYScDNm7O4sfd9WBRboyg3/7rMDPqvx+QwTBBUv0oxNJaQuNDfRzgqfg0iUypr40geQpnh1fbPy
Ct4KdFGcp/jDr3hsz5n5SwrHOlWWG2WK27IYjYIeuPIzU5/BPKw+sv523d8q921ATJWXr0Wlucfd
l+4Zj5jzpuGho77YpGiexCQ7Sod/KM2yJccKautYouneXfNnaVzwlZ4kWHcXEsbn+9rrwBSSPRWx
c73pKC3RQ6FezNV53nAeirVPt6AIJ0Yf4QxsOuOu2wuLr9afv5RdrBgQmdfUxNeRD74wQ/H2PxgW
SkL5Zb0hAxm6tZENvI1D4tl2I8ciCVf91OAeC1jZ/qgznpHDGj3un3ahbmGpCRo3YyJsVvm1rHt8
mSRA6dV0O7vi/IwqlvqkWrZgMxzOxfOvOEABGy0PdFDBhcaois2WnfDcnsa78ZctBiGoOnGg6Q9R
TkgdaSozIX446s6EfGm813EDSSm7BUDiKfwLmV0s8a6TyHxf0B+oZqGO6KdxZFFs3mu5nJ8JN4G1
l+JScqzMRV2PQIL+YPfm4bqDF9/x9zI38P3Qm1xCvh0w1EQTQAhy3cXi26b47TU3mGuXj967f7YY
9KP9TNEDNmK7Grayizh726yZhUBXNh5hZLYy7zsdV6KZpVFKyJZQ1Kc0GeSLjIUlZ/d2vJVILy+V
+Cfahd/Rs52hTmXwU5b1gGyctSlx+BMLVB+tIa73kdz1c8Mxe/ynzoqMVMkg2wQx7qsssdDvK0Ft
+qrUvvB/SD5/FwTW8aSmoUllWNgtSzs7Hihgm82V9x0Rqs2yWYzQ+LpbOPbi9+fbwdTuuI4+g3AY
W1Rdlw6y0fithrd6lHOqPf4oLV8VAF7ZQt1HdAzPFP2XB1zUh5SvggkXikiGXMgJ3t+wkGY8GXMF
JQrrWSJ0ZsXBRO9RuYahSmyjzMiHqaHFYB/bz0xg4JraiMEhQ76Hi8hJYyCEs0dh+zGQEP8xPTfF
yU50V64HTgINHnM6Vw8Brk5qzY8O/+ihXnYzt9hfjACFU9DRXMNnEZTwhApZrViSQ0ONUIrZnrCc
RN87VdWmY1HaAVqVuNOCszeipvhI64y5ngK4+ftRUkkCM5Ijbyy5YhN/GU42bpiEQJuyMz7GaRJy
U2siln/eE1AqU53S84DM9tJkU2KlwoOlAE/Qop5v3obOCnrHUZJrsEPX6Vnx9YjeePhMv/hF9drx
GLRO5RcZ0/V8PNmRPOjNKNysr9KIDLhVQ4zybNX1Xi2q3FhjzaKfsFps0DuRxV8nRdreaB5MFaaR
3Kl4zxlni7FORF9EiYweCuZgcp5A+/FNBMWAUvZtu8WasBkeexYGlSeBCGom0dzDj99AqcJwzXPL
FATj0/lMllHOU/5Ltml9yNnLsOivVVn6k5lSmfGsqkS9vWVBZFxiVzrevfufukGefFTc6Ba78slS
orcWL6lTH6gZnj56pnndhJQ38yfJ51663PXi5v1wMr/XNhe6Wb0sckagjDF4Lnah10TjW/J0Ctoz
5ahvDmpWSV8pVhtZt/Qwp/Z3Qw4JcHypFR7S6tJpn9S3Rch2KTK8qHsEZtMnU5bNEa3ELGB1vCuZ
BUp0bt3Wxpy6xRFgoQpNc9koDGHkYd7cFn5Kn9oVa48xDyNLyx8vHifRdR/N14CEtv7uYWKqn3Dw
odjvsUNE3NI1IOqZ/suOsv6alcpB/tAjr12luFzll+MzwoEQper664PMak+RqrDRiU6LhlGcJGy1
jc2xTj+1koq8mRTXsV2i3ofbrkrBpyBng6aMveuBXMS8tnXFlgsvaPD9i+d9pmYsK6WXfwy2zyoq
cD8sTVMWNbZOmwkBTRy7FhvEHT1d/mXGehkvNNS7G0ow0B2W8phEuZukIW9H6KAitt/GmOfJaUys
Gpp7Pa6CKAVn1FcrVjWm5jTZUxL93R/r2z0/xSgqN0RNRBuz09FmjLxtJl2MaC2FzQ6xRYWKWhJN
JWZyN9fA0sVWYTfWtLDhABFv1t+xFST4a09gkupsLHPy/8R+P7iaMjWPPEaAjID1s1Ou5XXEAPqY
E+qCyCLCo/1HKV5rkAM0wM05reQAMNiiE2oOzhSE7kIPnMkEN+bSWw83iAk01ZzDVHlqoXT/5p9+
FTzsKo8mO9rsfBaJbY8UUaYSs/09+x/kYPEVm4NV6TQ/53zi2iS4w6p5ga30eAbubV3Ekc5qQmsV
FmCZeD/zLdkU+YINKJLu/1XSf6/3IdbNMArtAUyhWudTe0IpIpM4e/fPl/cho3ycd5iemjveJFmG
tSX8BvI//0O1GI/XPYCRnpzWgoZPrh2A+ekpGarQwdID1tOf7zIGka5SRJ4md9G+FW0OLvVT3uO4
DpgD4NUWx4G8nZOuLp/cmZKdZTQoZc6vvmRXZlcGh4tOYJWx5ECtCqiUoZPhwe7ZEny2H5m1fVST
KN2OlNlrDZMCZLuuuEQir8987g92sn3/K4gofT9t+DcRDxwUBt6jhOSszXuMzP5iwNQNRGTicStj
iyiZOtM0qZabQRpTWswlzjfpKV1CEdVpgpTfZylBZfSK6mAbStBp2AAKeO68WT8EcRVHOY8SKmaU
0LqFKWup2jdUIsbs+HSwawgQTVwquUrjy84BEYLuxwngD7KS5lgrtWqA6ZvIMZ751XT88BIeO2lP
Rgo8wVvKgVm435VC/1sqqaEF1YqrX8LF3WXwhibijUC22Ywr5hjGapMygBnaIRCasxV+O7rDov8n
B1fzBP0FX1Zs14F2zi6ZtcfFovxq8MdhbTBqKvGtL8oKD3EXrXTNeukEuoeLUjZGMKPfwsCTPPjo
6fjq5whyM+ChwjFm5e1l9+P3WZoPqoK8+BL83PJCPfarbaR1rtTsOHbGKAk6SasYfgUPQlmrMdwb
XUMQGZ8JdWs4xQfG8liXFsI1P3z6p+Kiwxh15AjrUr1cHz9oEsvqaedD/UtggauPP44E0epo72NM
tRBEYPIqktJvPSXNl2CzQlJ/STtDwx/Obz3u7FvMFXX4BT6+FUKuKyReTWgZtdQJWTa+N7uB81n/
36smS9qsMByDetPqkBcBg9iBwhGsJatUqr+dl4Aw6dVe2nwTvtpcepv7bzkLaSQl83TkzTpeKL+F
F2umfjCrk2f9eSMdm2yCmvCbk5ZUQWDkvyB+bvddwgPsEKxZvj9AADUgmZjiiu9vlNLBm2xfKwi+
f21LICifHgxYqw0ftljWnd+lRkH9loQVJ8WmVkV5TuZgd2lH1Kd11j2bCJdj2qOI0IgfqL5jYeM1
5CCQ6DOjv/AafLKMEVz8qhD4RDnO8qkftOkA/ftB+IBLRnzYpfOu9kKi+9pvRmaGu2G11BPwyjr7
uoChRwPvQwLPL95s5Ju+6DWW8QWcLgzI6AJ1pXa2zavGkwbg9mDzX+HFUIywXn2ixnursN4lpmsZ
H5aYe5TalPfU5ieZHHHlAiqM9pGct1jlEsobcB53FKkB5zORCrir62lwU6xYJU5B6GjRzM47rY2L
2GZoRBfEdY0LH8n/FKhqMT4Bo0ooa9kgkFEVFSMDkbk0ZeZzUYav8cJTPbt/ULTPjVBLFg3MNb7q
xLTpNW82QJ1LoZy6NFfYAd2UmOkvqCxl41/DVtOfpQmFubQzH5vm6hAmHHX9V9gVPnh1IQuPSMVQ
WndFSFX3kFq9pqFZhu9kDM0rerartHw5NKfB2UM7dvQAvM3JeNL9RkthZbD0Mp6NXSJbKeNyCh7l
sD+FepJR3K+bYZlbij73bD5K6lkYK5LgI9C5DyO04bRh2jb9ATAec3dr8p9R6Vyyqne9pkjRmZiY
50JEzSwYnUimMS46W9+/zkDHvTY4ay0Wlx3jkpV8BsL52TJnWO0LB2A1w7FgBDHTcaxN54bTFhMH
tRln98X2xkqFpo5ggyil2ByM6mGw6q9phJ8beq0ao3/yrwlI49s3ag6UFBlEDiBkPkjhC7olssDr
gX2O3MF63BsCpww6a28lREaKhzj9dSml2rp8KmQz9xgFkQ+3EHI57CKczLTfO9ntHsFAEy2qjqIt
eFL5mvDHji/LeH18GG0E+drwu5wgs3D7fZoVNo0jcttbj510tdbAwc9+mQ3O86f0px+IT9TMPsbb
Bkmf/sgbIudXYKusrcmpg0kmrIWYInrUdo/HYSFKm8A3mKfr6xD4TXEuinHQi0EAF7/fbFelDn95
+97kEIp+EnxleqLztfWLGrd7j7FbB1sS+xa5ovkII7SaXCozIqn7OWVV4+FTYmnaJ094plorIcZE
E27k5IO4eu9LnoKn5rE6DRWU+EpMySjHO693HKPljyDuumLJpnl6UTiq/koghALCNCRmEH4WdTTO
os/REcn7j+fwNUiYsumYFNNh9ra2z76bZQfB4CLlkYIi0981ngfyoArjE+HMshSIG4qAw9oxfUD5
7XVzXgxjAQPIpkuIrv4RAoQmFU97dMuXJQgQIxe57jN3c5saLTUfhvT+UaqN8gB6Gn9gum8mlMQw
852DTb2lJXcY/5lC02kd+T4TrywLIoH/s38kR4hpDX6h9Egp7miSkkq05cfwp/LLrVHE1yLvUjiL
l7xRNxccnUhriLa2tLDcsqvNejuwoMZAhQ7I4/9Vcw6M9iAD3TMwneygFig6/B+EGPTG0QbwuXBW
Q5bd7W8e5A+wUWHba8X5AYp0Ys4Oq43zDOplxbTPqy2PLE8kbbWyESmzqFMz5aHX7oz2YEFtuGdw
FVj0Lnx+n5EGs56BkMzO6DXkUDZ1/txsqPI9f2+pbLEDBH1cGiYRaYwTSd0ItP9aS9nC0EGePDZn
fWuaJhiJ8WFL2FiIeRA8/0b4cysL8Sfjs6av+OJtYQRb6Ws06FFKORBT7PI79Keq+zaq/FRI+pRN
Yztr46ZctWCYiFN8e03Ujdo58NFv5/s/vLl8XDWZuLeoADsWI4sfGEtOPV0kJYjG6aKLq6nvOCTg
wsuR1S1XwZ4bVOAszgmutyar/3HFbFKYjmByADVqOg7FFjHybPjwIKzcUmaFfCz67cin2nS0gkg7
JR9e25NtGAAkS3VFsA3qYeMdGXTFDHYbqIlGLLDB33MMNuhBItGiFIhNzQtrpyDVfvKMvDek5fr3
aTzwQkW1lPBOiHJ+TZwvFQLeMj1P3q6Iw4Da8i1PoXPz05kubmTkU8P0I5stxPbhKvKXWZVgDdaj
pe75VqE4QRvpYsZumTbpIStqskLxZko59uG44mS5n/Vc4IMjqW3a4GAh+k+p7k9g0s81V+lNSjkD
FvnlTDsreHC2wB44okjoSOvujBwxxz68BbeD2Cz4UbwARwFwvpMaMCpN1rHpsboMuUei+J8LR3t9
ag7pEzkvAuZICUPpQMeQgFgM9SHDIj6wQQFuXupXzzTiXVkHjGwzeH3mCamHSQEnCVBQSvBWu2Si
3/eshUI1mwfX4ADlMvET3RPziYLF6FFovMgRnG9IywO8x8jXobBEJBvKwwksQUYT72QIw8bafIUT
pqY1dtS6SdJ/LxJp8Uw0A///H6Eg5ZGMafO635jMbPSxYmKvWiDpFDBn3djkiuZkvHNjaj61x3ey
4ePsF9n6ffTc4+qWf7fpKmyF2SG3bk4yy8DVRrIJ7tg/CMHMr/uf/25Qku+wBV3TSYnLejjxDgbX
53FomUdOJmAXWCsQqwliPhZMhy3bj1PH+ToZvy1NCQkwJ7ApY3YcvQvfXAovN6DISG2wo7NunZKw
r+QUN48RpY5ZVrtbgCPAMVSoCAArX9ozVJ5YTLYyO3cdzeg4mKegIu048CEYqx/wNQoysnkThRp2
Wlc3cJVq64ZdH/nYd78i3zVepvpixNEKeH5oy5YXQvKmQHUy3oOYPhkCPB5bjB+YuACPxUc5TKip
S6RELEPj1Ypb+EgZPMi7b+tfXxiFNYf0vdDNH36akAM4n3xBSP9AzM8UDxfXIQxdROpa+LL7ZH8+
4PvBe1dmNg3a8rar16lWCSI1bzh6MfpLZNXSUmLslQ5pEOhso9BwmtuT2t+Zc9daekQydQbjb5Gw
v1lcegG6RmvWNyG4+xRwJ+ZpO4zOWoXTYcq3IruAEsZPA9DxCFgVvOvMQS1BzG5zn3fyaZJte8gw
r/ts5/RJ3hN7T3bMk6Ij2v5mq1PxcIdFE+hpNuekzegEndOWzXKju0DgmxFktA86Hn0PnFGuAM7Q
hHbHY3xgA8WQqnwrtHK4bRsVl5E7ARjLRLi2qroeciwdwBj7OUJB/Iq9HGy1edbq5fwbtNwws1n0
NQiVvg44ox541hqeriwiW/rjpWzbHt5xbuMUjFbI+qjDzw+oGY9Pux+j+bkKnp3/zKJfKVoyKz3K
W0SKZ/2/Q+6Bo6Up6WZAKctbZWbvyO1Xph2DGj/+dCcEyMpigoaEWPlpWoSjOlgb2Z30MzSfc/0M
zrr/3ZuWdNjJIovRkFVMUIu9tlA8aLrfoqRL1eaJjREDX4nKpOACR+CV3sTg1y20bmPd5WB5CkSw
oK71V6vmm5FEyIFEYqmfKnG3CoIqY9CGyaJ0x1YLSFxDWvaw6mzUsC0HfshvfZc98l/Tf8sqotay
wBs5jk27AyN3psAqYIvFczy9NF3dFG+UM9qMbUtO8onTRjxX+eLlQL7oGp9/v89w+Vi+hHiBqYKL
YRjGRtcYEdeaUCV26rrtfxRyOvY5nGfK6dKkS0lnwrupGBA6EN9dscyI+LL7ch2VqUiiaJ2NTgSW
rv9Rvh928kW+AQo1yGSIp89nIK0NZivx2kuuof6tst39nET37/IhimtohkkTONpR7YQHT6VTW0ac
nwZ4d6isxc5iQb74lhmVOKZh6Hsi+rKVPNlJ7rWw+shlAydPC5sPj1c3D48UbsECk5qqj8/+ryXn
4bmD72ewF3H/pKRDrInB4d2yo/n5ljSiQm8frhfATGPOmn6+nh3fwOsI1aQLCxn5FBF58HQtNRbB
SGADqYosQ1p6FjxHP02UiwTP3VoWppRzWXZw5+3uI+pNmQbVsa82kyf0B4Np8cqgQ7xdDjrR2AML
rm/jPMWolm283wCxrsOfQwk3ThpBG87ilE8Etulkd467FoWqs8uOcukcn+pBT22FVrpuj0zsLVFQ
qUQ8IPU7k4RquOd+a7vCAR6OHvdZ/4yr4MppFGUHinyEkKw9V8U+aAnaFbSGaJBzVy+LTkY+MhrW
1h+Xg/o5rdBK9+pgof3ugFrvq76/cLdwveEiQo7Yq4mU6pkLtrDdQizt0OsUB84KjX11CSgiH79c
D+XfQGMmgDDR+MZgo6dAjsvVHPwheqTt7DRmodUPpiFXio5p/0tjEzQlco0+Kx59bsQ4ou37PaFj
4bTGDcwY1eJ1aIb5yLvtzO66C8Aa9Tag/JAgPIjCHxWFLx2foIOKweEar/rZ58+vf0wQPIbA3j55
7u2Vo3u1wnfXukg/lh+2oHfO9psHYOKxh8itYEs4LI1zNba3W+GKGPzLSe6wxA/Ma3cbUpefD/HT
WOqroZSU+LoxeqDDkU/YVvnI0UoL6CWebAyOp5JDGuwt2J9R4ivEHS5bVYhVJsQXn0BYfu1Ili/x
gdbq1ydnxwaIn4dEP0icEwHUeqZrtLa1YUxaxqN0V7OyHhYdZ6dSS64XCSBBsq53UkNWC53YLpNS
03bgv7cNfVPBdnsX9xXb2c+HsdLa9LvY/jADpWo2H00snC4IsFZe31N/D/mbNXealMDROXVM1G9C
IyY7rHdZNyYjqz60G2ipvcw+Fk1RTHZahpaZUPjJrXplCNmBFv1PZYIBeKqDRhKH3GSVu8EJ6jIH
LPWk7ruh6jOc7jBHyQ2kPfK3UCETj8CCrBWMM7Cc2sP8MHa/jDBEaGLQdzuHnbz8ir1pVnVmErK0
ohtZPj2LkHorS8P7gNc5O8Ce5WTaBmDXnd8HRBkdrWI15W7b+0n1ifN2kHgtcp2zgXH6GUmiig+5
ZpSAHYYIVt06scVoz0pWC+LOUH6ZCeFwJRb/ZOMnpYPFlLNWpk3GrrqMbD+43W4HsklZ1dC9i06Z
T5zsU27Bo+xawevzHGbi3xbWPt7JS9XK/am9RcodUKDxoWdJTDGrBn3mxKWkAJFVNrN0q/tPWnsS
ph4/fh6tDERNbqZwVCdtenGiFRQblboRZa9RosI3aAJcQBhOsrtkZSJ9mpQFVl1UkK3wC3Ik4MBq
mEx7E47wAPSiGmbeTFwa2dg7CJAy4mJJ8fus9HCPcsAo0TFgLVhlkBeVqGZFO2VVXHQs1Yssleyf
fTfShoPIAvY8yzxIFipHvhyts707Ku6Y97sYsxwnFqkL8z3EbiQvvcIScere88Vm/dtLshpRbJBp
v3MsWtRzFfpn/PeDjUYkA5BXNWBGs13b2RyVwu4kQvsmjNiMRK0+ikY6q0qYT+62/HWNmUKKe0lh
c8cLLPdKA9WahVLzOT7wEc5wFMDf5okDXvJyVssYm1I8gnSubcs0Y6wq5d91oha5tgTmEEiG+qWL
gCOey8BjwXXJKAkBk3MRCuwILVFYBWxHcatwaEriEKQY5JMzLUd+hVUDK4J1Eg8sKbU6qk1M01zQ
+JyAIRhlOyhar9POgAQGbSIIJjHiH6iaH6/fRXQpgBact561s241ea0DlebfXchpBOI8ovEQVJxm
7iA8uAw/oUe6MOcbVtFx7nCG3n0jVDKxh70AtEMV2LylLlb/26S1n2BAH6ippXrzQbxiufVzetvs
TFtijU7X6OcX2wuwoa10GDsmYzY+14YewPBitKswd/pzstOPMAh/nzBD61WtNEKyhZC3xq9oHS1t
FipveARoSTZtmydGNvoq2tsgfpcDQd8Y9MGLOp5OyWEcSdA4Qzn2Bfqx5Cqc2dzZ6aC6e4/RMFZ7
X6rILGs+d1yuXTjCWrfGne4IawBeTBPHBAg2jBv+qUR/Byj5MkBsa6tXfjga6ewkV2th/L1NIOPr
oFDb9OwmMdIIIg8B3XQ+4uVIU8xk8bT8ZxPj3CamZL977ZnlpvcpI204tWSrTCWaMNXkpdDSir3v
WinZUlhWIg24sNST6d4t2fY/4ymCv56ZzF8AzJZLo+J41TXdfSe2oF3EewTDqiphHMMkOgRo2LA4
Z3EGnLShK5EHcxEaHsVbS5iH7QKG29CTXBtxT8EVpgp7xg79Br1kNB8dLUq7qwPNBCPRI21BW10X
djEw2nOoj29p8pmi63wq/Jl/TZ1WmV4Vu8bXRKTYbbN8A3B6Uj1dyLayM8q1eGgRjGqYrCmZtT0K
dlEYCoEbEAwwCcdzweEsJgzdrcG5cDM9XQjFJDhvFtaA4i44VfaE487l3UnsWsFVRa7Ys67XF9xx
cYzfag6nYWKnwv9BKEUt1MEf1y2xs5em1Ist2Csz9C7y/VUMHMHBm1VZXrTdcthrm0G0bXtgmbTQ
resWnOX9/DwDB9GdqfqvmA93U9lFlFxC8+Q+SMMETF+MUGic7sK641wq6bA+5eMm4s09r4fkcyoz
Ii1ZlcnYtCaxHoSHjPee+Y/3FXxVbtGy7+mRJxa2EVxAIXlhZB516BKTMQ5hAGazSOhxSTW73XCS
mEvu0gp/7UmQWVugvk/bEfe/d3ktcyLiPCiFiWqvVkdabodt3kJHnBDP+nUMPKP6Iq0GxqnVFOa1
EnPPMCFqnAJVVMNBSegi4gjjQCXs4zDIIzUT7x9i9NakGqrUCA7xGandMq7+w5hbji2ryPWzwilJ
1WyC1SlrYXt8MmEgoIhqA011Oekwk9Ak9lXfSA+CrwwIFlv7+/FYTqJSmLyIWLgndA/HZ14v/0mn
dk5aD27J3cvPA34x9Ev5DP3v5vh7PI4JYNftP/Nl3rtTBaDT/vSk0HkqOlTj9a3NwqsQOOA9K/fE
qIe7Q25eFrWL6eJpTxuUcTkbyipRbL4+3+hP1bjUh+M/z1F//ZP3rw3+CZibvP7PZX85JsNpKwNa
GJLMrbIm6EsfOSX/7M7EraEeHp5t1HJVTWtLPHh2j5pN13gQzJRHdCOOIM9C35nzT8VQvMWa7Mtu
/tbYRSPxV+0lbPYZGQEvJu+vLa0sctNXbetE+h5lRKV0CS8rm1UvghUOfM/ZbkGMuo+CD83KZXQa
851XHAgzlgJ9ZIWZKiopm+gXKPPd1kAqgXnVxpSDAnIsNl2YQ8Zr87AOrWWDARaRMkRPYglWogJ6
htQtnB1aQzVSmpsJkuDEh+Ve4lQAgzlFtnNlDVLS6vBxtsl49FNc0dKlyH5jPLksrZ3V/tmqhbRZ
LTD1OuYRcVLjDPnNu/WAyGRnCXZvIKOr6Dy4aS9cBCgSklOBWxFNcBpAZbuAL96NP4hpyxcuMncO
K23zkX/kFStMG149YYLgveWvKQj3/+Gu/UWZWl1bA0e120KJqIpvKjhwcEskDHsrrzJAGnhw6SHi
090WL8mpeMWvnFZZRuyjDs/zVs/PnPdwNNBpCYYs/MiBQc+OyBjkyo+qCXsTZJjSVN/mAE8OgOpd
UYkZYLZB1JRG8KVBG/qMbSEawufwECYwYYs1Hgk3KowXWVgUa0NayI92o++XVySa94AckyyM2NCi
vJ4SYqqkACHYAyBMBiUeKprwrhp4CpVSYIgnNi1c5lTw3DxsGP9hw1bOrvs2AMaWJxvU9IOSLblf
JLY9SbxYeoKkzU0SdJSlIPmCiyGzazmE8U6Yxm5ICjTZ1ngIOhf72TEQ+ObQV8pyuAJnsvxhwbiF
Qn+N/US77fTB8gRch2/x6o5NtKuowlf6axMSK+BxtQgOzIlBAqVJH70oD8OV/1DoRr3CWbZDITzb
lQfTEvmhmRF57EuKhmb9wB2HvbSm9+92TTf+Cb7YAP+ziP2Zhb+VNOD0FkrE3DwHiEbk6StR0vYD
V2rOLT6+8UwTWjhSvTrME85PKTtXeD6/jznEhGO3HXdBO/7Fva7ph0N8A+9c3dQcG2bH6L0C4PXX
IJUADYJ0NLn9DoBFlUA3Nh01vkxnko+oRGWhKFcjLh0+rSYLp7N3KK9avWRVEad4kP5kQUFvIjsJ
awwHZO5tV4LHfS5Aiqf2OybLSk4IiO+kspOPYEbWQ18VfK50xE+0aZeLWQNwpzeaXTP6OFQ85aNO
MCz9vuES9RegvEArxGD18BP4m8XF/iy+9m4fXgnN3wQB2SnX98Jp06ztynemHLd/iYQh8QOVbGdE
V+t1rqXVu4Q7iXkTuTaKFZwNFBB6ziU4wqCSFhXNfJyDTIhgRVapts0f7fKKt9MOhUMh3hcRqywZ
Zoodj51WK+VDrZPmL9/Ux/Ifc2fxZ01BJUAqJxnQdpuVeQKGoWGxSLpjqRAZTvddopg968nCstuT
7S+mo1kFd986Xh5eBXKvQdiZWjdDqPvN68/MvO77xRyEPcPU+4D3DWKFEgZaMHPzfrkyV0/I+2RY
Gs9IMIDaW+NzA53SIHTsVoQIUMqSOME/xbDtVRI91qJcUy+03//N7xRNmgXt1jukvnVCByceCjTW
BTFGYtErLYVZ0AdtzVKBhIMglZWOPwCrI8Nm/CLLR3vqxOzaJOs+XyZ8F0A3TkZ7ov3aRE6pAYXm
b29kGfP/JN5z2xpdqmCDhNGivv2Q7ji7HwSkhDg3YDIuiDXrC3Lo/vQnx6OmmC9wabBwo6KkUdd3
K5kNekcQm47nLSfyFglelJBon/4zf9nm/EOs0f/Pb+T8SY7MP5Vei6qxhktqQQ7H7gKhrLk5muGd
qNRVET7LKp8GeLMeTi/CxfEMb+BBgENlV9wqmqrZ17FWFLQjoP19YkBGCOn2maITmJcR4JKkNSbD
n7AKSvkHGetgK6OOxIvtXQ/WegLVn083xYyvaa7qjO2GlWZFMqf4ad9WwSHvjmaA5H0GTsoHgFNX
Tg0B15a7RWGfpCStiagE1uNbYZP8QmLf1xC0Ozp1AnXHpXEABE80055AwrDBETzvCb1zPF1npB4t
Z7A51WNy18jsVJ7Bi5vHhkvO/xg1JRnYRuDmIJa2h0na3NKBBHr0UegGTLNukdx4Zk2/iEFVjBKE
gIMPFSZhvXmzHgXLPgCxMJKdqcQnW4DQ/KEUxvy/0V+V/CsltMi3v7X2XkRjwAI4ZJQUH4NCDzBm
n0BmM3qqfwJWBwy8DDwxfEaisu6LUyvkq/ZC3KN7N+1MZzG4W6/yv2fy1UTDbvHmiLHMxYn+FniD
FOZ9HLwHYiZPusw+1DV/Hpx5F0fXNuy3GIxWZqjqtGQlJt3tJUuOVIOQfDyHrKJJrFvpePGU+6MA
sq8s/mnqIek7i22RKNo2wlsfy6ZQydxcxAqjQAeKcTRMzp7QR+mN9D9L1YOPDXoQVnp3JQScHDgu
DcxJzR2Vksw4rlTn7vauN5v6vflm4hPMDK65tOZaMw0u9rCJBapesAnVQbgemMOs5f1yemUNdGH/
WFnnzbKSHJ8enXH408uMKaIZpSZPu0K6cX2R01+oOm2TsCtwEobVjUAyU5PsoAGGdwsYuTS/Qhzx
7OqDaTEVE6ojIbOdN5sOiJS2ItoEdPl7p79b0VhbPm2I1eb4RKvyf0pQFCl2NhNqs8JAExu4WNwD
iZS+w2+O7XumZZ/KH1UQ4+E752kMQX3HYrk1d4xQ+zwlS1c8G1nwboWig5xM4h9YzlZ4Nc+S6XQc
LbTpyZHgUIzuQFMYMWCrpcw9qQLEZJM/a/lYGGBJolHfFPcFwODdu3uUNoyBBpP6xH7U1YiWKOFI
BI2rl2seJq2fmFmhYQrvaKf6NZY0A+5BeHYGV40rfhX6CyWQo4PMtRt0Lxx0/WJDEkZ7q53m73XH
lT/fsU5EXWRKZJ6DXi3oV+uqhHEW6lzzFofKr1Ym7uo40JQwvVscGT82lFC5b9Jnp8t35FWhqnFo
s7d4TtX6pC+809IW27cppW34KCCdxiYfQBPgUxSU3b3vfxLTzed+eJKAR9hhCJbVqj/Za+lfBgEu
OEwwmgFeAkeSlx+oqT9cUeaJ4ndzoXbGeORMM0Fxb9OganchDTbiCQ9c852SbrPZGcbRdMBcvTnU
e2SQVlOhptneTXe1QgTZUU+sjrj6LyRxS1nVWybQ8wXCKG23dkVYdpKbgYZFZd9anfN9AEI8gCdb
AqMrr67uly+RgiRm8L069FlOksNSsfZOyn848JVzfaZXg3hvqIs9IwQs4aZTPxDS8MH6j8k59Skq
dyx9N1WobCi43P8MUqlsJGk0pdoZCPddiXQVjlCSgHw9EW9qYXnjVEmcVmbVg9Ab4XPNz5aIfwSM
ZtsKnK/Ah3wbHCa+jjHljwwtoLb1aeriXnm9vMcX3NrRnOtD5kGpHBAdBFHM3lQxqM0x1qoRxZSf
Rc861ECKgW5QFns5EDb766ABq1WyrTTkAF5adRl+o+GR7mkw1AZ0UB+WODcUyy5dqLoTY8ymHH/+
LlI8H+2O5czXO/kAJeBMTQWSD8peNfAlCY4LRe34po7LSND1qFL38b/oi12yRaYmJA9ir4GwzqcG
ESSH8h9dwQ/VHs1XmzE5XMLB4h87UMcfS9/JuxF6Om5G+sJBZpYmpb8O+3XXR/MUgqVRuLOXPXBi
u0/cxRSHIukwN+ycHbvnBhsfR3hy4Xwje12z1ejCIY/oJPUxgshHsGkXQDCRk4anESm7A2szpUbd
jT99u/9mJfFTOy1BWIUPHO9aZQv43sJ1G9FvtzddlqJ6J0eVC8EboMMNM1iBE5zp+Dg5oPCSKg7N
joVrYyzp0YILO2I3aIsOefchyUZkX5XfBF57BY5eQEhfSStWFjCoXqhaXeoudrYSb4cBNdnoznVe
dZS/4K7uhACWEwN50Ek+0whkb3uLOYBw7n+W3GhSAi+w/+QjwbtvO3JLGBvvJb8uKvFsuXFmc18n
BgpLQT2LsoV+3oxJTj6sHL5LVaPDJodzN+4roHEpyzdPND1tHh6MDCdlrsOQArzGxtP2KNG4/MBR
uIM7WKOkKNvoatShsJlMsvL3ZFPWol/csHozXjcRUO2wuPrlC/yuptqv78YSG/x97Fl0xdPDFXss
PArO/Q3/SJWmZqRNThLyREvfpU2E8kKF6csVt3UosUb7/8lSKYdRexOCa/Ayu1B5qN+OrXJW8M5r
1+hdfm9y6Br2fpbNVrIr9ha4dWZ0pSGZF7t3yuimDAUoxHfLnPSWtHfsZN5gEGMhcZ808x011MNp
4cK/ngZRjt8xpsBoxYRwWxs8EObAyd33JSSuOmrH95+tNWsPydHG8vKvSaEBoJlNVWaVr9jMiR1d
FNKs5bBg/MAk7mSdDv2v/DG5D2GfeofegxL3gW85/dmT707RVH5xugz3BPpYqcE3Y6fQI0MKoU5s
CglTr9cHHUM7Rp+on6X6NSc2o3CsWsNMp2wp8e00tswI3p/DBjjfOWoZmxf6ddO9F6PLwabvrBTx
EIDkor6fXnqy5G3dsy77MGA6oTDPuwl5g82OnbAyEmssjNPx41NwGPrnHRNtJsStltkOh+TAHwGI
EbQ8Qhtr5Zbs+IdHuT7h8ZBCjLyp/E0XY2QZY1FwPk0Sy2GDaTWyJCvoSCQ4BOCY3eU9Mgjt2cHf
fZ01QWPpMhurs4zYNGMmixigTMAjCifonkIVLiMUHqaPIHaExfNfiMmyY3vhjT7JhNDzVDFkKkQx
cVnkf7Qe/bth50XCaiauFT+8puGz7e4DIiHGTEs653y3zUgINbrduNVZswKUsDedo/i26/rtGATT
p6d6Bq3ziLRFhFwruX/83tKr48JTg+4Cuckxrg+rSng1nxs07knvAerlmejptGwnopMBBzE4sMZ0
HHx+8j11F4LHgrepwvB+FXmx1qw5CSkc5upgekcWjjkc6a4sWoakqemHflAcR1BYCmNecZrzuGiL
omvSy1TxHcqvAn+yKCX1bJc8yc0/Mce2ozjcjhWOMaK8tZ3G5SA0at5GO67a2x0LjZatFTa17cNi
L6BToNZJN4YmJgaufghxjCUZ/xXdpaL0qLJbGZ+xp3TuTYz5ehSwlG0NQ7iqFjnAJqjpJSM2lQwL
j6og7TqUJR8vOuxRPOTaYOJZiRWz9q5H9FZVcoJl5kXFaxFl/mM/4y0TtBvHJfGivoa/Z5xpbbcM
oDPgQry5EJ1FKO0+8DGSQwVPu7Usgau3wtCIBnw2cTkX3ZXcmbIXJowCSYsveNpBkMFEVbI8ekvL
rU9PcAiSWp85rrf6KsX3ZhpAf6xsDV0qJ8ECAmfOv3eDhyENHJZzF1kOYnzGJjzUbwiUiUoKfZxa
8UzAHyF0zqnYQiGSFzbrcCMSK2cG76Q7l4U2wuMRpFGgbR3fYE3GjJC+fscC2HBkFL1HY6jAsgg2
NSHEHZRYEPUoshsn0DxIDC3nIpSZqMUE3HesYKfwuo3wtvyfktF2yc51c8FnbMv6f4Wt+nl55UHY
fAX/gUXc70P7IFBKXwi+DgPKTw2oMnftpuvVqI/afXTetjo5/YkaHAciFCdgkLP8K6hNWknrdaq6
t+CeYrWspXdz8blq3ZlEHAs2ntHyKgxSoWY/6J9ESrBUJk06XoPoDG8iP/FSjzQ5Oc3Jv+Ipxpci
UUigNyXrA7pYwjmMZnJbVB9Q+5mA46/vJzW4Ch241P+vzHQ4qaAhppBKGPQjTbLGOkqONWcy5VIl
LJSvgujY/1CDh+OL5duxa5cW6P8nOjPCxE6huwt65/ZD6+kPkHR1yp42FeXztvA8hgYUd/YIG4I/
5PhgtmAs8yk+O8lqwQ8qvNL6bnCISNIhRRrI8ibAhUXWmET23xdmNOouY8KGlI/Jy2gF1/aULeko
vc3s+ATVN+ZwuHRt0+Lf7SSY6uRLA7zbz/fu064DG/fXvfZA9PLoJrsqv2rnVDBKE88ZQhqLP6ND
F+1axY+F2PexMXkhQFIJo7BFornCx32W8ZCRYg/b7jb8CAx6oCPHUGdeeDnXyRr5MWUr71+h7XQF
6xbojx5ceocscQv02E4aAzBFFj7K58hJEwct80zdCD6VAUHRKttnJObN5UpgjJl0ZYnLu6hzNjEy
Xj7NO6LyIXgoOYX5vOlFV91oPSAzjailmL+d9pnGU8f6qdiK+nNvEzSr/7aVLOjMN2nVY5eN1i/K
BWlJEqInS1u2N3D5d9ZI89IJwPVP9yeVuijPKGIgywEsME26d2b2Qht/d9iOLQ4MsoHZTlluyBy3
D5xUZayE8w+MHImGcObNt4tXvw9/R5uCDItgZP/m9g1szo/QrAjP3dsZ24HaQTKP3W6MdHt1LN5e
K+9mo+Ofs2+I3mG/RROT3qW3zbgBpM1YkYxwMnBKsx9oQaNkXqOAz6X8yzkXtbFXwNYRUKnwvZGG
W+MRMIsGrqIurH4u72Q+MHaln3ysWrKsZn8P8CDNlOKLbuWWZUJVcjs/C6U4VT/HsnKlaQEJU2L9
gGedf6w3uYAs1Ktp2xBxPt8JlobTzfznmgotbjC8JhdSJY1j/m1TL7hsWun2D3yTP4SfXnn50/Wl
sKMD27EXpEI5KRrVspBwOLhUI3qkRXi37pNg4c9oJvACkfym1+OiZkePEka16IhT8bMzlMThnUgY
ssY5Fc6E4dPjz1DYlQ2oqANAoiQWsygv2RQpj5lca/IFZoOjBgBj9Yd7h/uV4Ev22MyptM9HTG75
zDNA7asyH22+xoWbztPCfYYtqdAZqOqKz0nVHhC5EkdYoQE6wbsNhODyFNL7Dp+InC2cAzHyAxPK
qr1Vrb1IyjOeGDY59f/vcN1QtoIlbcumtL1YcVaMWuRBYpufyylH35a6zXA8Ow77EmXwO7lRzx7n
4sBcSgyuq6j/n8gHkxqUTweCUTigZDPPLYvk5wPghfL7jvrc+hnZ0TQjoq0oV/8ewtKwqVJXuFmW
q3Wg3m8PaHrrkamBDozXn9cFSZEseD/0fsxBm/TyzTFIFJJ6vXOXadgcWCYNBieodWBvqIvbzYyN
Z/QMJkFKgW6Avhkc4MRuoatgwdwILhbJbU4EtbBiC2NQ5x4hHGd+IxvXAM9w+8Ci8FmIH//s7v6v
UruWl6FKQD3xL1PQzEIHP+Y5c5z8XayS+qPjLEuPQai1tUmppgc27RcxefQtfGQk20pSE8ld0TXq
tbkKkAxMCnTXHVhswLR0V+zKr/23Xc6nYkYzFLkqb+sNpqExGQvyC3tqjc8XiDnCc4NC2d3q4TL1
4rrXkmVnnh5WGHzvDXb9fScmYn47z48kdbd9WlT2um9DpF++GvweKyii8g+NKpUXbDu/QhKD7NRG
74P8VlCq3+KXMruIPglizB8X7coNbmps7PwenlLG54CVQfq5FsbzBZr/QI9D6oW1+lABXd74UZmj
Df1ldFoXtMBaxKH7d1ww8UY3VNohm2oW4tEPYu5LnwI46iBViPWZ0ApFkpz9LF3h68ECphwXOx25
iCgKvEyhmBKLZfYPnwFfPs191XgkmYyTVlhoWZGylAJYzLkGkMQ+U8LLy13Q7/WYHsmznF30T22b
XGZw2v6v3NgN0wWUdi6B8S5TKCpYPwdckK/KrSqJi2UGnWLf7dxb7WoZW7jY6WaPXkjpSlwMr32/
C2gwbiEoewQ+OvJwGTuODhQFw6LKQYO3ZjL8gdZHNva9SB+TqJg0VvgzHJW7tUoxLmWKJhrhc4Xs
mIGfTudJrsfvWasXO5WUxsqOtTGQiHvCaHZaNiz1mfxaXEcSioM2eElKf43w4cfMrpJqUEIf6FCy
ZaZ1+9UVDDxcufdKVp2Pps8tK3M6OEnkMIRz656kas5HDn3GfT4/N7x1Ne8i1e2029IlDJGffNXT
JPvrqord4DPyeMrSADbo5bEeEK29LsQtmHH+E5cEDmL667IWCD8fYap2hCmb8/+CRLGHh9KGsxYi
Qpsnhyy2KO4h8IL68jn1u+8F/By3cmbPW7juf1fbuyzvHf6Lp4T4Ii87IMx/o7Ev/QCO5Uy6zAA6
g8k5MHJ8jFUJvt7Q4FVFJwj2Pig7+OH8Ffxhybp8ZKPw9zosvEXaYMnSXHh6RPBoU8sVV0wtBoAQ
kGEt2hrDsVeUojkkiSVM6HjNkKUcqLsOaT212BxTaO+eVbsXQbb5FXs7amrmRWWoG7t257zestyi
3KOWYyZ/Tyidrdm5G4y1frDw8ygTJe4tOWm+opL0ElZMAob1jABGov0gkMFRLcrJ20/fABYGDmSt
JteYlrglhz65jY8UO6Au6c9f9upnba/NwdGu31XMub8hn3kmc/VLJLnhW6VsxUCcs+vdm9yEL+kl
R/mclHeh1afbvn+NEPeATHQIUDgsWq7MhgV7mjGTG/tam2tXxkz0Qr0LZ8aKonKusT//wNN+zKMY
kGj/W5dFnbftJgBYvuMu7F3egwkGesOy1DGD3gnWrMM4DbCFZwR37ts5m3Yebr2PXyRdyaIDw4xZ
uRHlfbIbqqeFQJjrhzEsos/b4NavrPy+/NbNnQR8/VgUbwVcbr4ZKOcCb9UNC0mSMvz95OWQUbEY
T0CSUz0JcxDvOPPbR87KSKGzQiyswQyqkiBxnToMiJRdzEpgMomKlobb11P3m5MjOHKV37kC3B6k
KAvYpAZ2I4kBGXLqCV3zEpbiSI5ARBYuF93NQ2hd7El7nVpelmSujj6mW3M/+GvcBJzNGnZfp89t
Py9u1T4PQy1d2Qu6en1M0MKyKin6xeD+Jhz6PvWEpLviVOe24yZRMMXU96Vu28W7/kHyAlXNAYEk
HTGrQH9esOQ2w1wZ19lCbvPtUEBw+FPdkwI7OM+wxasKrom1ADYC/Stfw7uWESM1nSayAg/2K7fC
VwFphV+qflnsHgPAhLW5oGbfJx/xTDh91NLaL7KRKrEs7xkwuROdJtDGPBAAtc3+6dGO0OUGPv/3
77PUxVp618uJA0JS9pW8aj2NJxPRFOlv7tWCnRTswD0Pdb6lrT7/ev2zNxSm2Flcryer7+YXHpQJ
kr+vPI2AhgtoUbCUGg+Tpb84TJcuSkn1tt/zu+duZ678LSYbXjI5VG6dlcRQJ11e7aKbg/0LOl6F
D2jeVdgXg2x4ss0XjS/GKYpziImwqj8fKjN4REHMPTn7Ce1UmFrERn3b3/K4Zq9g32rJ18cHRw5u
BUSxVwBDvYqfmstonfFxCMddIaqRDB9rwEhHEUDZDMTNcLisASft5rQdm0+Xp1YfT7syMqKeIpKC
R2crFCrrsmZK4aLQylDIkFmvMiTshsYkh4GMEIc6wPJVrAcg6DFx6X/WyoMD7T9YZubaWHunalGi
fqHcqc8dNaUADbjD+FvFYvUqLdHhOQph+5+nmRciAYyslZ5opzOSZFqwJ7uGcKoranMoKvCF39Hf
i2rHb94G6B06c2/MyVpXbT5HG+g5gvWyesIXRGVD36pBPC4wzldDS3GG0Oa5AJL3Zj/pmHlSJB96
fg4jVUp9TlN+S/hXDQ4c3jujGSzwfjJd/vZl3dGE1XABtxC0+aQ7Hl61zlDawoUHsF2XomezVx9h
wf3lWDWyfmubmRMEHFNrX6Mq5bqSlFkbpZ5aSantag2ff0hpYZWe8DoTJj+Tx+4gDBBIkZgFncgE
7QLpocccEvtHlEzJQFKEsnpF7j09qsC3GDQmiR3j7ClTn8cCMXzzxESkKoewCvhfGg6MDnwjuQdH
d7kfgnLmZu5Iq89GcPB8BaUSB8SEdqaWj/8rhwBA4A1MOiJ+ZIVbe5W8zewKASIdo9UZ6IF1o36Y
DEIOMAyBwiP+L98/txJgs37hGOnP6NXPmTL33IsaTkApHZRQfCmw2PIFoHOQLSSd83D7IIk9D7vx
ag8TlB8rnwuhNWvk/OUl1vztyK+jkDcFStSorqK+RodCIBgm5eulNAxHxerGhUlcj8fdHBaV/9A/
7xySivGhuhZjkygdFeHM2kvIVj7vBikDU434bIOuMv30Jvtum1XAeoZStb3Bf4eH+fR5+YEjc+li
mr8RvZA/rYMdU3dknZoLdPMkgR9mahe5RV52Q6NdNHU4V30buiNk5gagDhGwsyAMfZiookGcxhZs
6Sz9H/ImAjaUE5USV5tMxcuxsAns+H/S9zjiSwDz2diISrgQ82i3zDp789Jww0mEkvTjktq4h+5m
3lwePS7enPdQvVGJ/Jp2ZYVffaIqUo/lx147Qhv17Wmd2Kf7lPAbPDNOUOItImTtVUGzC8pxi7XW
gSRQhCWQelicVOCNRJ/PFwX4obUXSq/5+f8ETdikg+hssjqKf6qe4HHmYTNmsEWgkQlh7btKcVC3
21q6fwlLW3kcce8pVMikhofpnKfbrg+/6c9ub2oKnnOG6mBfO/ra3o4K99UDbo2hupWarg7+aHPC
qwNkV6VXxRLGBs8XIJ2G/jMNXhX6rTEcu4tFJ03EPSCx2GgzFHcWufGRNDnV26NZhudJff3ZyiA8
4alsMM23d+iNmKabTA4cxiDORWR+sy/xM6mEbwRXlOcMkQqlAN8Vr1aO9i5+wPqd+u8dN7HeJ3wh
KeiJxTS0KvSt/dHY3cKCFPhcs0q6DxYtlU53F3xVCZFGcFRCTe058iLtm2kBEabdx5x4ltHXoH63
bRAhP8p2G+pc8c3fTq5Z8igdA6cWvya7ZjWquy7Tnu7/VO6rKBvnRKm/ZILYDXjupMAmOpjlbyX0
nfrvY6Cse5dnp/a9f/1RL5V4zo4xBW8d98YKzHDFAN0uBi/BDlMAVS04WK2lNgFoyiB9yxeUMv1R
AzalsUW4GBU/OE39fHg36MZfU50V2zWDet5UV0IaL+Mq3fc12AD6PgXZFXfUidNlfxZADa+7DLmz
Nd51mztxWx70HHIAfs0cBF7/SZ+Z2iKJ6qDWxsYwtnBkOYamK4EiMExQeaOcvWHaHshFA9mTL1TF
NHDZ2qNchDtOmg4T2z/eFQ34aPr8FY0nciQRBuN1zhEx1Mu7aE9J1LcA+wb5+MhRNCOx1JOsioZC
jNxrhMGRT+z0pE0AAY9iaECABXkaBe1vIi6nvEmGgP9Wgt8dkDnkAEwVbNicpqCKk0t1brs1yxH/
lqp/AlPWPDTMNw1GbQG0LCEPHFFPqMNAOAmuu/p+1NpXdNBdlCyU4TwQM2tSFfOTGbILu3fOm3zK
bDMgiCPU45iUkl0HEDXRKb6/WXxpa5Ml/VPUPu/djIiKuLmZWlpq0JbuBdrljLy7Mug2iEhvkPOv
9lN5g4wnc8Mp0WBJJR6vhmMP9flb1dMJKuqWPmT3eL7Sr/G1s+xorf0SFSL5H4HrkhZESIXuRFDV
6GMAc7RnnekVdxkmHLbnMPOvT30dSX1rCfky8hT4yJC3IbTJX3R/jqBz2QUjFazHotzpQt+uScU7
ZHrX09Xv58IoGtJjZaXER5Hapt1SI7T5CgdCkCZawvaorBc3XYqCvg8yNrB7ec0K172Ai2d2y9XP
xH/eW6+5NrSHxcsC8Ppme+/2PS2PU8EwM7J9VdFda1jC5KCQ4xg4T1eyY10B/mA0WYgrt+2gOL40
3Bf8Rsm2uT/wMbV1OpLDycfl9UPMO0C4MuOF7wa7uNLir5CSUzeZwsYx4bVlf8X2CqMf2UnrkhRX
nSoW4MD4rE8icqyJrIc3k6o22F4dWony4n/+kK8lungNf4aCbewP6LtnJh7HMF1ISlvku9VTWnsK
gFD7m2Isfk20QHp4HvkRBOkDyCVurkXZzw4CAhhkjLr2TQ2xh+2rk7YdGeDiUZtRjVduGZeEym4q
nSK+1YF6Dxpnio9ig6O77u6owRTTilZ8/S4MQPK7r14tPW3HNstSkWHIeABpxK4FtWMRhUlswdxQ
ru0wnLDqZ5IDsFU7/dXlkEBr0vYeBK3O+xM35XeF0vx6gldg5AJkt3fz8P1ry3E028hWvTkQyGqL
amG5beNb1tTiBvLhochXed06T38P+23INtKFXprbtWldMPHgfTCYr5oyqJy2Rm/k24lP0mi3IYvI
wa1OTa4QVMtkgTNnVZpz0oSSpbLQs8SFcLF8x/u3LmAg/xz0rbEq3A78U66f5+A9k3lCUQyIQLSw
m4okJu8/GSPB6P6aIopn8/EZPpWpI4xLYm9nRTO4R+o22nybZA4V2F8N9itZp9u1Ps31GRGMcoOc
O50ex/+6rWHD+1PHv6VK+TY26z2yvzI9zG0Rj69GzwMrDUS8oJq0ahELQN9zTLOl2Xv0TUEGSINy
9plsv/KI8jC+SK2uWkl4IWCvyHri2UWUDiSbjEX9Bcder8PmZyDgpdNYrWJJ1vVkyIXUftonMQ65
L2BJo+jj/SW6rMFsKbGmWNDhzXoaZin5D6NXi1BzIzD2aDyBdinRAT8r5w2eibfE6zNBFVOsamQN
lEc/OBHgc/B0BYXZi0C1TczCOtXHwRpjTe7XVpSH3SDqcs9GGfb1C6SHVM7FL98/x8+Osrt8gQHw
TRKgCiiEZfufi0DtVMSgRewsiUjbTPgfFoxAPaOzBlExUJFkMCALiYsChx4sF4lTMXznQqxVM56K
CtP1elYBWZm6hwAux3ecPah0ZnD6RkwApSt36jB5zR9nqEDkUXtma3mJYqTLkAbzxZecwWhqXnei
34ntfhLyjxDF8wUOkssHZq18/5JtQ54N/poomgGKY5/9hT5Uf23obg5/cNu6xz3yM7nrCoKzf++n
u9UfLH5j8sQN68N3s10vQ2vFeeD6/HiH/e25I67AY78teaZ74wf7oJjEYh4JqDEHEOcw4VCWEvzL
HWfNftMx/Z1NfXL8P+MJ/6bNdBI8qEwfidlz88vhu9IDslcIlbYsah5JU0nCkz+C9Y0obR1rpefK
iWfZ8Po+QniFMUtuRBbSmhZiVhCPcI5YtmW5pD4oVN+zkFxeD1XNvUDGg5Nu81gpG2D16B5bYL9r
m1m5Nd+xBE5sHeCFHm6a2Vgi7DK7H9R3pybUyp1/l58RSXFE6WGGvfMQeFo0g0oX2RMp6YA7biwC
kFfWCBHeUWU+RLXYiWjysVADegXOIkTD0IbBJTOnoWVchGB98MjDyIqRdcXYEL3d/7lnsRsvejxp
lRCxqiPR711tTzMmQwAMsgmB4YMfNDgm/18cpxltjw0vIYqtU5/7dDjiVimZccHZaJYd6yAkPU5a
A1ME8HMq+oLQsZcCOZL/jWRyNoAptz5+uip2rZB7roktWkgyQjdCyuSTWjpFPAJZP952uLl1ypcz
rXFaY+2hpLp8lZqgjnqIpjBkaB5zzaEMcd7gUINE6Ss4eh2LakZwo2HSVzzGTezVqZPDD3w7AGhu
QDCAM8yF2/dQYNjX2oiGfYJu/CammL1Ft5jvufNKHGCUaGxpdXEmVfKuVPQyh7ldP14CZCQGjISm
MDVbu9+0sKsFFmddTUriJW6fK3+n818Z2dHGYO4J2SGX9CVPDi5/J2fnZ2oYz8Gc8cCJSAQJNUx2
pgvPNsO8pJogJZNTrEY0eTWpUf8b8CnTneoAdoj3uKpslV+i7LL8cM/HWJroiDYCkvScoT6tXgqn
vUz66RRh61ULcrvo6+np6VoLozirkDceIEPjTCBZK3Ho0JO780Yhti2Vhm5WLlIpfP4u6ZSqWuZl
YUGW1SIRQMjADzKtAKhC3YGpryDHXKa0kGl9XLNgcAhWNwtxZez1hfCkeLSfAf8IYOnS6wS8LFsy
dtJcBDJhFvqnAbD3FjiVyQCjcBqjgPa4jv6ODkhubm0zctVDumw8tPgylvWUTSPhvQ/pj0BZ9Bo8
TSzyaHOgOVWIKM8q3a3p27x7Gpt1tW1VSG118i8HH0ofoQd6ThnB/D3M+BhpCPZN0dGZ/e/7gnLt
Dv5s02M8l3Ng1a+1oQNVTGjdDfvniiuv8H2KLA1aWdU3am3uNMWVelRedL+HE9/7Xdw88KjfcIoM
SNjh+eZdKsiAEXSgyhvIfifR/nXM1/o4ZCQiRkNr6QvEo2X2bQDFPv5AhxzhRB7Zf1A82fzdYVNU
8upCo7XXsJpZ2Hx0By7L4KvrU1ynAd0w+fbcUBn1uKf1PeAUK9rOlWTeSws5Fjyk63jMCC1/fKzA
Vi21uNlcYwZqP7tf8V4HabAMia9QwlY6lGOAXOB8LDc84orf+9FwrmhYkAQr47o4JzgYd5RM55OT
IC+JOwLb6wuBfB/+XdCgIQUiDMv7MKHH6TLSlbxn3OsHPxW5KnVxOMJUFAUkDkAAVuJvVrPj5aTU
dnC+AeL9wnMwRi2xVRlSrk1WOdEvC7p4/yWv3xSv8YHNemceiGUU08CkHDzrsdLrOkdsh49u42hV
iWfmL/np0iTI/00xcNbP0EM85Nn6KHZxz3LE4Xo76ICG9N1OAu3XRzdOKw3fq3axNAPffwNFeMaA
Q+XZUQ/dulNXQ6RkL9Y1Hws3Nx2+ixp432jHZG46JefB+zf5TA0+c6eRdzkbjsD2b+Q7W0psH7ap
vu73IzfK8YIYoabt36rOVTmM0QlE82QrWi46GKgN4wWWz2k4/1R93JnFFvAsOiqg1Sh8OrVoByjF
g8e61Ocew2gyxXxZInbiejtWuCWI/wZhsk7fviP52ZCv4R74bb3FYugbYPH8hV//yuiumneB/yv6
g3ehLOkksMPawK2zZyMaqZRx8lg1QyshjWsVR1hxUEq7FyxpywDlnK3vU6uUzWyXppqqqEoprhgK
bHKp4mmXLMoh+gZcnKb9xFjgByHiu97CBr4M5FVUdcQrOzy+ukEN/DOmGw4JL43Fl6GkhQaUSRlp
MXtPp75fTVA2RUO7SSkyPN1le0onHGBn6feBlhgMz8MZnKiYfln/kA8Sacjd00ldRLdD6gv+ZdM+
tJVg2w5VK10MBFssmE0Fb5PNtjj6NCOWll6mPGykrp18KemgKIaVxpplGkcqQ+CKzSZ0hfNTArzO
dE8GwKiBNQN/Dr2ld+Mi9DsOAU6PGMIpJcnc4Z5PYr2cbEwhssGPVl2Obj7ml8/0scTAVxhh2TOC
JcXGudm6pzM+iUlWLSytgmW0HfRvP9vVVqywUFJ1oVf618LxN5uLSY3OZoSn+tPUMdi+7+ifAn6/
kNinOEEk8O+QGt3eM3bPcvpw6YPrU8SRRal+iVJ7ipMOcFPjuqmOoTiSTOl12yZ6ayZDFh5oUTNz
C1T5gCNbObvQeydXm3w9/2iPKKCv214BXeWNHbPm8BN/y6CRRpEMw/5PlMRh5E/zTDtvP49azGzv
eGKyzKndfsihUXQeETWLX0nTEPEgd+m1wpw/hgp6+U/VTOVDP6KXsGi2wV1Q9d9K5/nqfCRM0qpl
zhUq7OrLByWCDFQXyEqokWN4JgMvnUp5ELR5EUo1k4NePzcqhsLhM9ITLmq9qFsyYtWzfYlIE/WL
nUe/V2+6JZ+Np4oHaqXXtgnRJZBl9eydvUtFuudhq7ZL46YJvk9DKW2u2fFsgyepkus3vsf1NCIG
UyIdb6RVK2Zh+NoyW3Y0p3EPbNmem4pSLMd9kFczoBt2oT2wfEr6yBkuvIWUxYqFfc16x8uLEHwf
VFikRHO1ew/IqXwbwcZ0UTp1XXdKZPZV0W8WL3KmlkC6Vqh8leigglFO/P5o8FsIuvI873FXPWy1
/aUeUOA5DA36ZKOdLrYbVr0BAdr9vMzSFzZqe/F47H3eBRt8opHn/FOGwUEVF6MT4vwwwKclRqlH
Fttff2g1cOo5o0neP3X93J6LrlWHE0G0WJB1gqBC8sjPGINopz+34PIYQwiOdKr6Xjx+XuyKnbE2
+XlPz/SPWYD2o+NBpivP+mhUR4ysmwPHF85x6OC3L513HjLOns1xMaUSzyBA7WqL6b1FOV9pcavQ
lH7PYC2Pa93scNOIiQpSkE9X0qXWsBjVHQSma/c+qb+oUi3RT96VZy2mtHmK1j59USqGHKWGCkT8
eNnuL4MZI7aaw8itDybR9ocx1siJPHU/W3di3vWQbmpnTRzQZ/V8218hfasQPXJLgNclrp4splMx
YMvZNtI5Ob5cN9+8yzQfnje3FQVeUmI5KeKerCXaCqOtuuF6rSItxGEHk0En8JYQyQXsckZcoYt5
176AXP6UpLsYAVyxg2TNMpM5X/gfWIwGZlXuiLEyZV3o3EsnaMcCMXc7WjDyfhyW3oaX/fzKWIC9
EwrQikXPHKPqpFlbTwkaZb+oW9gagcEBQH0eja3uRtieq6if5NRwdT4mW5u4xaonUCeUqAPwS7YS
W5qGBCpl7rADwoJiY+FZPxh5vIfz7fpHAxTeQc700MjSJhHPYHlDFa5v32uf1PegUioU7vtBI5z/
bD+aD+dS0oMSkA8LbFSnOGJPbmuykU7uCtiitKl8yZGZ423ByXh07WPgZvRWbO2OxUvfdwUZw824
96WgeGDg47UYSw9QHWNhR/sHXl9c4drNlttHswOd9CKCnjhamOEKQgpFWQ81B7IH+oI7JRsp2UHX
wS2Vqyekj9FKWiKQU7btzUpaOdfQZbAS2bMCEQhIUF/H49dl1NYnJWKCLLaaC/h3CzYkKfNFHRwJ
0wUzRfspltRYC1dS0Zk6jsEmiA/MSFUBOqyvTGJj1xiCtRXqQR6nBnOvAPmR2FMK9dVDoLalQ5fc
M4WDL0Cx2OTVfH2fgt8gBy6wedJVDYyH3zE5LSq6H2o/VxkCDCN6w0dXZwCiyC3+71M+z7ayyeCF
qOAltRmcNWmCUMEcDjbpm33uLkwiYuI0pJaoGcTC+2qLZnxnsBAJIs+PVuknfr8hPuQXLTtUyf+6
z5wdb7vXLtkCXU2dGnak/iPHgwk24DIZRinGehdnM9ThxgfnCX6Y341D2SOvu5RqgJzXde5U5Zxc
jYSZOWEKL+oo70zpIskIkEBH+9LOYACMVtmfeNOgroBuw9p4vxwYwNiC30S+G85zxjXpoi/gPV5h
jTNL0VPWxVZHapoUtqF4AYtK0n3nBOJzTPwm9ZRl8dh0gse7W3wSVOqmfEJxyqJm+iY9/HpQ957/
a259D6pUPskBc30ckvNqKM4AqtmxZNr77dCe2wMJsC57ig/xqfsHSs5uMXuINj0Qmcql1HvNThJh
WqQbJJtHKZPqq0w2Xfyj6dIhI52TDV2oONtSU198wODUfGdLH2oVkoqaYuWuhrPi8uL3BsatUMKq
LJUeujzjNZw92lXfZliO6/k4AMtNojNqQ7mRbmx5Nu3+QiQNSD5JW9Zs0XaW5UUvBayF+FaAMsVF
9k5TEfEQ/5iGgakjAn+MJqBQECvuD+cxiCZ6Ehyy2armhm9vMKknH7yKxISXkRkQcvGIaTHuju6k
CbUsuzH8vYZozVG4F9l8sm5iaxRrwYAkaILdbLiu+OhThAxboY05g2CKiuouSCc6uJjmrISnwk6E
w/hMzvdN64jByTp6kOI+/mRtOTwd+icuO3R2s0LZYsXFA4vPnm9+rTAl5mroMaDcGFA1D6noOaWH
iU9IocpX2FIcGqUnV/SVnV6kMyQ6cMA8bBRo75xq9mADe1gawURtCJFyzZAUt0dj04rhSOtTo2CC
iPnB5am0qllFK4ADhQ8aueveanZwnXFt7x9QZblg1AvPAOBW7DtW0KlL/Cx1i6JBlYa3cNsWQK2M
whxYQzxu8p43Fy4zObVlMfo7RUNjUIf82ToTygfMDADOpftnbH/s+lWEeQpCFTE7hel+7kZUns+a
aeEFUKG2yI7RnhgnniPbevqtmRfdZfewDIg/upGaqzC8UX3PWCb1swfCRWn9Hx4bHR58OZ/IgJwW
noAAbEOmK6mTPTOBN2d84GQd0d+B7rgjmIv8tVFqygiED4P84kkFnLadTqdXJf6TK5/fUtBXmWqR
NMAuSGyw4hwHBEy7/fDOxWyIsRAucjUV3UqzuuaFJ8m9AUgFFHwHiarRClYQ7NsBakT2jPwJ+ECR
kQGZEP6Dm6jCD1Ws+rjh1VLloRQhsiPFszdsYDKoYUAc8RwzZ1UQayrXf/E7pNfkcNmMel61DQB3
uIp4XutrMYXm0wNW9I0fwzUGIlhmIP8f8yljV1XCy8/Q/C1Z2u+FWTK6jIe2FsL+Y5X/Sh+fXzud
fSrfLtmALcJU81BimG/AQMwJlROt92juHtLMiUrI6QJI/1AQbhz87y0+1SPf1UmU1pUEEfOgl405
rD09bKTqKwd3JwtVnoraurL3imK32iB48H87gBk1Do2x7k6oXpDliTcODvqBHKLxo/FwCjbRlkYl
/bKw8R90kRDgpv7H8A6vB9PWsGXNDCRXVWoOeUJwObVCI/X5hWMgBwbyc0vmIrb244cATp9/ofdi
KwYrBpO1un50p2lqSroi7YkcuU1hD9djB4+YcSxEOkLTTT0fjqXh4FXTqtR3X0Ft8jaF30ZuKa3O
YbjCJikAEse5yJSIIFc0MtQEgs/RsoNAmW9wclGUxvkaM7OEIWYDUSGwYmqazdrORdF/dJ5i5B9B
c0obhCRvWNgHWzdBGWDqDKTRzNx+SQfh2kaU4SlD9JIighQtLOeVGiL+jDiSsO+m34unUtHEETGm
9ifN9BHbIkO7mUxJk3dOjW6ZS+pONO2sTsbny5wzJu1bQnwFckRSg0RqmuVygfxw9Wwn8wiqm2bh
vA34JVYdCO/kHTVLMlHuhxNxv/77WOd7u4VRPLTiF2SRzZz+JNZfWihbNA50CnLtrqOTxIwgji7l
h9q63SdsntZ/tVkNsSRw+CYPvQ1LPZkbrH9rt9u28rP3yX0m6NqFXZ7LvGCB2lN7e7dKINR8k+1p
Chcf8l5XMsWW3dtF8yJefB0fR13Ks0awKkSfXLQ+QwSCHw9hqJ/QdfkoKPVGzpo+0DPZW4IDP6F1
+734Dp6jU/L3FqR8JG+V+D5aAu8/wHiEDM6BvzS8wyoEO+8O7ZnhnMWHyidp3TXdh56y4o/YRl0L
2c4JriyI7n2RLwm2iCfNuAHcO8V7D8Hw6nbzw2m3BLMrxKa1YQ96LU1pg7YOGKBb/kjrlOCZCtN+
pYXA/ZRXjNc+pf7SZzD2KGHuTQFB5+NxHfL2ROsx2vOG61Pn6fSj6Ev07z84yZGsvgBa+nyA9a1C
lvwuykF7YQvfniN7ROzBNexPfhAFJ6kaQLeAcxCLXMfZPsW1XHu6GDrg7W8qRt1lyClvMnRTwZGk
TEnoRBpvrxLUsCTDiKER2XjVZ3vg4C9Wxwl3YfewFCjRkRv44PQWbA2mzOPE/DxgmbbZ9u+/s3Zx
/rHvHSGrqSh+A3KaEobCvVRrlAxgnDxkpVsqBKNSygETL1FRMd4BKUoxrx057BAIu+EqmWBr1ymi
+LG4mC2sRdeyh3je0KlfI389ZRV6frfj9udLBsIvMLuL7CQBxKIp1EBA8Roztdp/HjkuDFINKdJU
nNFjbVVPqlHJVB79vpRPbDKiIyts0LsI7osDFTzOgY35VsMPcKkbUF1hYO7IPm1Gv44nCJitaOlz
lmZG8e7xtx+bGPNOrz/ZdV0y7Gz+ksTYg9zckd+GW41OPiI0KotzJOaEQndk57Am2lYBMwT1Y/Kr
HEYSY6KZqCEBDJy30+Tz4hVw9PUgKjV0ZfDIGt8fFPEOsWgpdv6iLjPT0Zw/67pPUcSE5g33UvTC
47nKk4gKaHnw/Svh1FM2fG+EgS3f+CNRnS7tbeb8rmv63j7Y02HSNJzdEAO4UqP9nlmx1R/U5iGT
QQehHOJpZlN3UehEbv73Zwipkvc+s/g3h8vwaaWOYoupB6WmQVOSkw4o7CP7brXMdcDpJkpT3hBm
bmNO12qc0c2WbMO6/Nwn8DrI3IalyPvfo+t4iUv30BpOZL4purIYQPII4eghL1+IGVwgJNTZgZAC
yC0yjaIJAJQZRoZF26ZKXssGJFCFht9nNs/cVPE5T2Pxq1zdU5otAbFrzRawZex0UI+0ZdKmKv1+
oi5AgChbPtnWPrRMxzXmi7ICEkx7SeRjIPEejM/kqNh7xiwbKgXZ0Jzq0BFagb1Dj/UOvH441Gtf
7p+EGAaOljuEW3h5WudLh8Ha7uUB1rnaRr+LbUdBtYZIHuu9l2Olw4f1+uEGHKgH9trSLvjPyfGw
OhGJ43i8ix1MZct7TyodT+1Dix8c6Al1tO/0wO6b0RDU3sYD3QzoiyiSwL3kh7CPriWCyu9ysmOb
4rxe+wT2GTq+kY4SpX+R+4eZMgePW1rbWnO156BaShAdTKN6Iip+VtoG5knnpYbP2wv16tMBsIX6
qLYn2kEIwAcy8ZYYTBtFWXZwEQfRmixsgp+7RRYtTY4Gx+devjBya4IBAB2bWMtHj+kL4Ktzt7Zz
5xGKL2t8iJ1dwTLv4WeSL5trpGeOpt3N1FumPVH/wNz0AY216YCgoHjby6zHLVOiZzYxrlQ3XC34
qjmbMCCTguCTej/UCW2eJgS+lmcZdW1Mk9wOfWcXJrG86bFwX9tAEp1CEFaqXCkPUoWAVugZJ80G
fR/su150H5AwhmCL5QxuxgeRuOPQvWJiIerDU4yEPNjM1oY7KKTuZyNxGIO9mierRmZulevmTMI0
VdoWSjb+4FGH0tu2RZtFvWpvzgvQ/PgaJ1vF2DvXDeSweqivnk4xjyiC0REcQuD1KJnzKn7AyNg4
mG2kbw7TvokDlu+kBsMnzu/qufncGuscqiYYBukxdgd9dDGX26s7wuyUDFqoH4wIrUbuuD2zTXdZ
4g6pqE1g7xz4wGOWJfaBh3D/zGF9b9dL12JAu1e5rIppcowpcht82cQZa+Suq9dK+wC4xwOc+k8D
YcOLLTdP8xJ0BEsrByWZnokDIi1ICgIoKet+n/kDlvfPDrwCRBgUSvkspaqnhF6KvS4nD2vQyib8
rBE/H/UunSXI5JfQG1FseO93h1mETJLXHJHgIbFg1gbxOVEU1hOqkBuH7ljshvQ759iBUfTn2728
aqIPBWmWxiaowuKAn55evA1EB8iEoBQcoqFdUkeQiewpctq2Bgz9uh9QLVIghxleluOImXmVnLoX
9uHFci/BBxke2lGujzVA1QbtJZx02VxhQCeYPkfmOtxAc96VIV07XZak24i+sNoPd3GLjwoloA+9
TFB1ajbJlyI0qNeoICps4+BgKTekMSkzKu6jgJSrSuFcOcTsKiBFf5R+u0um7NqyNz6I9QFMpuk+
T8c7aNpiPxKMhDyawHYMwyXDtYaLtM+N9rvdJsPL7j7BugZkV6CNHNnYoEXvynWQ+jg4IxDb1F8x
K9aQJzhsv+m2zjEYfMj4jFilDtwIO7egFMQxdFCTFgROaphalwyyB+2ftDKS14szVI1nfMxnRaP+
ozSjjFL9xt8cxzrzXWMHUINRNgcRyzgOeOkxKeY+yo/kMTHBoL9yr0fnYrT+wkITvaiGofwJQNdx
Rm1x6uFACJuPhTrSdwPn8EKg/aR8LwU46dxuKDKdy295StCbPG4iVLJVaXtHiPZmmbIfKuvl0dTh
jCJ9AJJIHCia07k+OGLzmi2sWMQRtqYs7yuwJPg/gM2kqLb5Kp5F0p0RN2AIEhU8hqmYQ2jrgGfl
6mWUEZZit73DedPlMX5/nlFY1fMhzn98t85QJGV0UjNC/a5ykO/RAOZ+NBP2LQxnRdOpbYPOSr1j
hrggsUEVHwUaNawNgqOcqztkETXJ4JN7QYI34Pl4gkvvHG6hJip8lKlDBwoTXIr8WOMvPuo4Ugc1
atDgYKB7Sq2hlpx+8+ZWn4k8kvtsPv1K9JsG0nqeZDyhmt1rm+uJzco5MIYz7MAeX1r0/Bn9xfyJ
p10+j+2xfIX4gvHuRrV/xl48ffvwUEnCX7iAbXTy0thbRcFqXZkKHc76Mb3ZKXoiFiIKCmHT6Pt9
3HcsOQS+Ar1QHJvEDRMlhLS5u9rgifV5KwPN+vz41Fae8LgF51ZPUbIUytgB3IRMBNefZCrbnWVF
n95EwGmmF8sYpB7BbGu782sSfsDQ9MTub307vq2lByvqsDLsJY7CO6vFtyUACgq6xw5i1MCgZ8Sz
Cw3ZEMfX1GJ9h1NLcU5hZjiuwk9TPeYQjneYK1oYabMm9W6kMzcTnPcoyhG97WdTBDYX+sfr0M7n
RBT2KnYZDKAdB9MZyF4U/iP0iB4yoBIgN5R9QUwO+daINhvRwdmqSB7AHvdlqSzIwoGUKQ8BE8e0
PfxnOUcULKxHxI0tX00Q7d8bfECYZxUOnMzClMzCKiglt5z+rD4czHUonzw2p6nO1YgdhJu3hrWA
V0wZqG0QYGXtFQhEpmfnL+K+aVvDfmjWar1fCFP8MIGeH2/QW/2NfBcAm63VRtaoVOtuxm6HwBNG
wLBpgFD9SSSQtRYCuUsrG/gis2GlfsyviREn1Jna94zmDByhrpoYLkHEyAX94aoPK5uO5Fq0K/GQ
lT0B6Eng2pjPsa/YHV/vUEa3g0DFncGN1aU3PGPA1RV9jbpcucV7n2pjz9PVSB3dNqMtTt/bo+25
40UN+VNip84pdBJ9UG1aeuCOrBR/8KcYbuQFT03UBShEgJZoV57lvAigv81LOoIPb9kKpLM8b9or
83jKphLZka2iVaZUIZmWS1BD1YRZ49Yx26Zhaq92Oy1PbIqVvd5CTve60WvwC5SByAm4nQLYUuzv
3sVUPWxliW6HG1BXsL3Akx5GE2Ngcd+5B0nGvg9XHZPOEvZ9EEQeIA8Y8Jc1gINEpRADCtxviL0h
hGN1a/czqbf57ucKiR5etN5Zz02VzRypTWgDH0tmhhb0pd1QNXHXjRfKwmHypy0GzzQUbnDf65E5
vljWL8XhlAswyE4OcGQ2phZYk0LH7x8AiFLfLO37jziedMcnfnJZLWNv8akESvmisszmRvLip7au
bvXlYCpPD7VbGH3Pe6rzpB7cXHIsr1txU19TbA3vp423f8LgEp5TANSzpoG3Zh1v/TUXrTZzvTfr
hznlEkmg6piieryRTZgQNtroSjv1xof26Tvg0lfFUowQ0p8KQv1xT1RU+nMWGSUQ2E69vPGZz99y
qWo7s53mL32Wu0MpkXbES88QSiNREBi5m40vAWIPIHZSK9jRsKZzd4wX3AxxT7tT8cWCcj2w8x2b
AZLgi3sz50dwgv+N5mhr8vuDq6Tde8At6f7+S4TAm4o2bn7C3VC2CO8IgMIqyRPLib3U0/Rv4D7U
7JTFOGykYkDQtn1BsfAfkbYmHy5D2izcJmhXj9Sh9l9pI5gz6YQL+chGkeL3woO0QzmffdE5fk+k
gSyYXz5H48cyCdLzhf4S+Nl2WZVd43ZEokXidYmNDVi3aMfgUGjtKBJtxaCdUyI0cp+a9NdI8Y9M
xTy9VOixoQsyr9rCjZ4ALCdckt8qFy7YeGyi7L0BHhwVAyL+chdoaYg9uHjstnFgp28LUwd6SKqw
4tBwnsp9gVx9qyXODCB8/uk2F2WAQLVxDbGtFm4X14C8NLVmU8lZiHjXtCeGer/u7S1R44C0rbig
Vzaojq1b9eNnkSLtrtB4xe4FgUCuV+mqQ3hZf9YqdTS6jS/oARcVScmqGFRQiFyYrnPwsbS1ohqQ
Tk/O9eoPK01mIopscjqd7aY1L/3IS6XZImnFAZJK+of9Yfls+0YJA1P2Qz7amvWSa28RMsSHOBkR
GMEeHPjgKJFr1wplDp453AKwu6lqb8D4SxwT1b1oJLA3/Qn0qEOugnh8ngOx1X+t/9ecpnJaK9s3
9YjpJJ8+QQ9XFXLDD4upwUlWd55ToDN0eL33fSRVXziON5FfUEHEtV+QPYVuMjojpboAJFIDPVGa
/zx5fWyE9xymONTE5UIx4Dc32ueiwxznLxX/N6WBn/0wKUUORALALNcCzRDHzE7IazCDB/406VOm
HdRhmgBNUu36MB6VooinBM83iqE8LrP08iF81v8EpyPkIaAYyksLJHgs8PYopE8MfH6XdO1TLKqR
VLP05kW7ONIj+9fM+SwfR07MUoljjVQf6HLxixUhPmVgSxZBMN1tK0ro8KETwiA5k7e0N39OxAjW
3mk+P+8NuG7z20sBOliI3YeNSbbfCJ6owWMsDqCBM1VPocG9ApuA5GHBG7dwLGt0ZSAf7yGZv/RE
c2DZqQ+/GOeoWjQHNSkWXqpHd7q3Mmi6yVLCIUhlzidI/zPGUTcG+UEAwl79OTDRLisbGELjOQu3
4c+IR053uaYqWWEczEXQF/q40h1VwBAg8BAHTHIFJ6hJfcMr/POs9tT+1pnWoI7InmPOcQpxKgZ0
F1QEuTSSipJHG7FeD/g3kQZLEQvxZA8p9JDqG2mnwmTt2UQrfehLqgQobE2ZwmBjLuTfwZl4/vCU
9WNqWYAo1Do2t18abbM44SrcGUqAzTj6naj9AGFEbZLHs/FxDePpJkBvtNJUZ3TRrH8Syka+siKn
o8WZrbFdUZV5vJ9HBxg+KaC7DJaVcDg5Xq14Zii4igHEbMutwSf2/SatTt6qDSwZC4nKMBSLeYaR
Q7nB4i8MWRVtyPmN5qBJtJDoJhQCXWjHhPZfpxJE1UzDiDOBp8a28CDlVlrk/hWjFtRtTNWSabfu
ABA/E29VU2DBnXFoDqWKJzwfuJw+JfCIk42d6IFv9tESKAqbUzWQpTdYvJbtIekz75rJCeWZsbFm
GQ2EWwIdYlHLB8+3ypcqWEo04yOZ/hBBeiCqN9tSC02MRyFh8qMgemjdke17dEzjkRbNXPzcp4jH
1fI7CDXcus8GdDIJFjWCD0NLwzbmadR27arldF0eWruzMF6ncemZWtWSKaqlrhoqS7J2Ko6qLmtl
iuEGnDP9c1nvfxRowjX+lhFGPwJ/WKOJmdQIzAnCMExZxd5tCQualOlr55S8XGosQUTXYvS3W9vs
J1ZNb9FATGGXIG/O4puAE5XlP7UEraAUy9OdtETQB10zXEEyuhbSDO2+CFY0gqoZ3ZAWAWvOuv3n
tOsYgTe9OOaDAwgeT/buIo3LG348Sfl36Vx198DUMfy/WExOwiWMHPgCO4sAVZt7ZHoxJh+qZpuz
OdHgVUKgHGCGyYuwP/11jAd7A/Br9vUYPnkY0wQiZ3Wb2uzWBSuHvaylNqiMBW0/BP3ieWaeYnwg
rZYxBwqwuczMIm0SqtD4qC0WO3smOcilcmotjF4CwfsnvHx1+k28NMVFWfb4A4J2zu0eUHNZtu9s
GaCQsdBm+/8X5XjIti//FcGbadmGKK455RQ6dVFCA9jwJox8paBeB9vzejjOPyRBUnmTIwlcmEuU
yR8yP8XuVZWlrB4Wgp21YT4n+7xdN6pdsgNZBqnRdUB1fNGrDuh1zff/ASl3QHUtWl1jxmEmyyuV
T4DYwzunri2Om661C3NqGb+S1QhVggz1EGm0zOxtlLqKu7ryPBhDOq+1OditAiqdGW92PJjOqLU2
3gfV1N+MPXCeqEAoWBIik1ExMwavujknhjxsIhOwUvsjtGkTEdIgIAlYLCa3/VSO29FjrbAXHBcy
6BeEAyEiLWF0H+gMu7jUmqukEV/9O9MXIgJfdmGlJn7oGoucBTKtlkIrjLvyURBTcRs8mSVHMMOl
P9cxgQNTby0QVpkyzsO7Qo4j47gKsmI6eVjUfqOWJ8f7zwY7touUWbwd8iNHbYHclZzrkh1Up7zm
nBNyrOeuobiH85jHsp/c0OhJD8UCZkblxh/C/DKVHT7euBJmFukkYfUdcYG3lcJo4xqylwbP1vAF
wmHFGrTazY6XrZvBOL1Pu0a5cmp0Is/Gij5NHPMx5+W2NBav5Y1FYiUXkHPUem9mj6rdcSD84wcO
mkh4C2JQnMpA8ZTxfQqu/Fv9c+G9nkQqAtqxy5v29CiK9DHmUQUKS958yYZHYBbZsXPq7P/F2vdP
qAJ1O+R4ZM3zjjc1FXo8YlTGiD/YH+ND5+t5oIXLBMbR3rDk7P+hRJ1jPRJb2ptXmiD8gvJDMt98
034l/B5TycmAekl+a40B2G3xab/FQYlyd/XBKBixkxGgeOBJZHnPBzeQue/I67gInn+B7l0VNtaK
M22AjDN//E2gsYDwAeiYGZAT7BbZKPW5omFmfXtaoVOUqQRI3wPE/ED1rj1mw9GOlO1AwVjZnjU6
8CI1nX7cHjxW0zJkPBneaclXzG7vyBKmcTP6T83ZUmAMytj2hWEegT5gGqCMtimUM8sSyJ5uvxK8
Qk6QLwIdOTI6l2lnFv4pLiYv0H2n6dNjlv75JBY0xvGRSqvSkOUCAEeo6OKVvZZfgoSAZm9GdWUe
qKIOKSjDixbxXKMlEKJyg+BVHby25UiWqbHNt8gNU2KKEGBXlHfEzgoAEAwkevOSt+V93cf36WZ4
H2/2zkS32SMlVG203fe7Jf68LWCin47aBkeS68dNmv9M30J8t5FET/i5ce+fz98QAbXI2dsbaJAf
JIr/Wb7pYBeL4NGx5uBs1xrzMdF/7OpDPFiFPCrS85qgqYGkuIlgWnbhBbIR9gtCM2hPSqZWbW6S
o5DdNiL/KJOSbm2wAx5k+yNjWcGdJ646gwWawN7bFPTzJnco1kmNzyIy8b4vlPZ+gLzWBARqFAGu
HvvQnb00qKnE3J+Fkx611S3tUteg35zU4/vtFffmKoX1CqswcPwyGNGgr7DBilCiodwXyNlj3thJ
f31BiWDZ8Vdq1wPVM8w52Z97YziWn72PbHfe4xmQcMBB/cZ5pQW7PZQGcoxa77+MD5AApygihcXH
L+AGsu43U9XzHmKmYinAxAQC9rYHf0I5iNzAKXc2YXp2ITdo49TaSlcNI6nyd9VC7lw1iVzrGQRy
4Z3U2fZ3v8159f/rtQ+NppRnO0G2sBsT9sCYHMwNNddkBqguuoOt7UVu2dozK7gyljUN8WAlhD26
QfyzHv6tDUKGSD3mNUIaf+O4jfGQPkPhunD2wZ2TuJlh0Hj2+dtlszdGXRBMgpfL35zXaGNDZjB7
4D+apFjRHBlgAEHpf2a0eRJwPROU2sZArKF2fS/Yi7Z5U2dgmOqodVTVSElrEO0F27Xx1zsZmyAd
YPM2eS4pw8Us4/v5oiHOyStJWmBHN+hwZlAJsji13cuEahWtPL6pvlKkNixGhcq25p8aW5uSjVbn
i15wO9tzw+JAPZg1jQ+il0seULuhNwTgm1Dpt+3sC/XxA4pMrEerGnfhbABhS2j2WYPKVyFXNA6s
jYbM4mzOadQtqCckoFZEc8UX+EU52c/L+Os3gNqq4eU/gYn1VC6h8mZMcu3q6Xyt2vWyVbfhGVEk
mzVob1uUC3lizFPGcsmw4vapl628XC23nJia0tz6kVJjQt+aKS3bwdZjc1iBm30eGeDlljs42me0
B0LMxlEJ3OJDYGWDKv5mg98TZnaS3N5ZqOLWvxeoJPFPcdkHODOsX876ec2z09o0xNiok10le0+C
FclgnkHDcC+R2Xb+6HJc5yH5OeRmlVrPWV/y6t88CClhtr1+/w+mxaLxJf8hCC4Yv7ZAUVmyZibL
CO9s9RLsOWEBUJUioWt1XUjAz/QQizB4YXt4vsmWFyzTrPdpFcfhINNFG5LaPXtsZ3l8+rwN4+aU
MiMs3jurunH9oTXsMSHhaHWPNNYGlBKs/qPeNAQLp/EeeqtV+JR8/RFx4Qh6PbNqzcv+Hhvr4nx+
7Juk47oTTu9QY8QBKYFuE3nBtMgU4fFuTWSTCuPLzqXysFAmMjY0UeWhWJ0jWmyIBrPAcoLm3FUm
z+AzpaRPPYWR3cH1vXOCA20P44sewAhl6wzGSpuc4B1hv4Q+5Q2BYxbY45TLTJKFU7RTz0XtoCh6
Nf2l3aoimhjyOv6GCWOYyNZZue9XTeauvj5NxlqugIj8bHglDfOR61GQgrHKFRmfZWrnNuJgrNHF
74DnfE5D4H+FIS0mD/thTOX92Anp/oieZtqSTyPGPLz+bUdgOsxUzu0dMFnN8jWpE99AxEQ74Baw
mucb65rlfqnroIwdQEY9uhCXF+iUoLj1pycxiieNvOpQUX/fTSKDwSpLUZPvBzKdof1TZOnj1qh1
r+gDaab4G2JRa9gcAEhxkS7g40NwX5H+Lblk78whgP7mGD+lru6NOfBzzmGzz1z87DiYfibIQxXy
ipDN4kPt5Bf38Tt6XAnHE5nEAPyiiLDl3/qkpotPYl2OkGOC6rot08DKhxYVfc+xJDOzPqS4osyI
n3Oha0snxFusKNNOtQCP36gkNacb2IzpTsJeVm6WMyuiXUjC19KGDxPR4nJFzLKytzvRVLspQNx9
LYiD/HhAe9L7vHkDkolVg/3sHzpCg2M1tbYblwfVnVMDfY2t2jHQ/JDEnOJxA3HLFWq4y3NLob5a
95sQnUyMoZIuDp+0kRhoSWXGUeUGafUTrobyFrFtLBAN45e9WepmnXGMPBvo5gXriVr97x3z3sZn
tGclolQcWsob/c3xIPyxVrBW2OXrwdwBEDyBm683Ane/0InFocV4r2vZt5Iw/MGchaIGe3N/t635
S6NqGMhyL1IHCiFUB/PufdLCx0IisWnfumB9uXM3Vp2BXLtc7w2fCJ+hXZgLUPRiJlxIWBy/bnJb
aR7+eE3Rp/VwOFyFYifw4E+0US083MTv7+WGLwVzd8coQ+xn28ETmV6o0os5wrfrfHprqpSOnIgD
63LxIotIeMBkCCWdfXTLQCLs3eX724+FsrOPFaHMxS1UwMGf7XvzBOKZEato1bnIxU/vGN1QvfWa
+OOhcpCdyoYUIl7ipJvOlgzmIYoNbfucIqaZa4VfMphEAQ1D5FfFwKqOxqjrg7d0+l8PzubGiFHT
A5z1oxFOYfxF4rivGhPrs1iuI6t1pLAJ6UoNBKrxhPUhUJuQkRqIppf4oh5ln1VW03tvE0+oMF9k
sk4b2AOIkRmeWKFwvGNaV+5+AAdSkRXK/47y4dZZLD8BsxrhPRsdX/P7dai4CSTn5OwnkrZ75/F0
NTAbKlswpZz/Z6zOkVOehMCbdlXSB/1smyxj9X+UlRHzBZ3TK15gyAtJ7rOMVMTN74HrS6WUQom7
huB1jrUE75gDgEBpgrTOvu0gmBycxjdlU2+oA6zHk6wgfP9DfovvrAHnHsEw8TIVUzCg04HWEo2K
nckqO20BmHmp54WOnHdhnmLiTW00Chr/LaPKiLScR2v4SXnM0YcmditBXHimIm2UB1vVR71FtFT/
l0A1GXuDBsYdj8s5BQ92SR4eh7SkmQ52TuBeAt/AN/pbs+FSUijmg8a1bqy2TcpfZJcaPel4Efjg
ZRLiTeIOmWTQJ/DKEgG8h9Hrvk4Mz4A4H4KQejO2/8PQs5eob0zlP9Vedrehke0ynvHmpIaqy/Qi
v5atF4FQKo0567Alt8ta9+/4IkOszhRwknn8zgAgcqniUSW8fD9nFD4oRNCCFodp5H1MJV1TwvH8
rSZIkQ/MatIWr9Fy7FBQwRGvQMqlPL1Q2DiY8y8LNtoJ0C8dmML3jA3J0aHZTdEnTA2L1vcibHvN
u/8eFF62CGo3P8rh6NJH6MnvARiZ95yP5smOopLuQKGsmBDakVN17gPd8UL5jyLX/7kDMRY1ceNb
VfuLpVklVG4wzjBm76z2IL6qCDsranZwXOnNg45qPweU+wiRoPtHN7VFnhjTzhtstlA5/3sD/Vvp
Ll/sAIqlaEOl3sqRXLEHmZz3xBRiMrQgAg+mQRuQFoVMALDZtU462CvY4QzzeZNrGhdf0H6XlQ+d
KbmHYCIQpBXoq5KSmbXTxP8G4sbIQG8n4rWW5x7rV9MFICqaDM81YwFi/D0GCnewrJmls/eMbZ+5
z+2tHzvNP0OAQugA+s5c4nGhJtrfmL7kimY2/7XQzc44LS3JXr5ew9K9Usa2K80hJkZ4NERsS+Os
eFL/CYKqFq6Hk0bNN4w1eTxhesC1wZJOUvIygpJSKc5EoFWMqLMYj1L4CKn8XTiiuNGZmpzBmQ1J
jw6y9AWwK2TiRoX1pBmYzg42VL7UQh9t58QQpHLgTzwSjH7OuXgyWKkA7TJKO7JgiCeMGMMcf2ty
6vqZWU5uHatb3YTCQHygdojBmcZA6rWgIKsQrSgJU6TLqUmLJ0apI//akXQ8o0EnT0kayemscGBh
uX8NN1wz+AVAv7Q5htNW/8dhVddotmGPxMfx/Cq3OMp/o3jcXLW1Ju2I0YESte58e7UE/5SV8WFY
mfZUGUmVpLlnewp84cXMFWsB+poR79JJAzOaXhv5igfPmq13wOO/ZlW2m1ueU5Xr4JuJXPtoiTcD
dZDV9TfMRQc7Elf3EulH/p5CwcslOmFRMPw7i2fkQmgbhDaD/aKeMUv6QZ9aTg4Q09cEyi7ur0l0
mkswRK0xbduEmrnhO5git3dawgbQkeguqpmLSPKhaSohF0NeumZikoT/JWTgn5U1XTgzK3mddoIP
rdM8d/5/JI8DL7IjWbS/ccBiYU5s3eM/kqQ3Wk4TZ0GGQxbSJXffZdLyI9I17TI6akF0jH62Z2gi
tJPAdKPj2Pu+5A/63f0shzpI1WDYIl2NE6VmA74pouOpiSdCrbbTRSgAUxyGQI7hKyHtDgR/naYf
KBkxFXoOp/fCiMdawR33t7haBZ1bZO3wZZSkiOm9DjpZ8K41YKZOteGxJYMChc6uRJv8wCcwFPt0
H6SwypcBcrXztQqObjPaqKQ9XM/DGC191GL+qTrXpap4s+BHKLNuQZ+xaZvwj4wN0HYfQU2UoqIN
PfSHdLrunkOaGlXDpHh+vz+f04ZZNpJYEwHlF+T+g/K5Um/3GKD3wGzExbGXhYgUtAwlZU6TWyy+
wkvWAvPi/JFnokG1rvwEkbmHXofZJy2ISI3plIqEA8+HI/A3QRqV01XUu+WCZJ1uSEOOKAuFS8x0
eEPucASmGw46OD04Fq3SVvVGwzagZ+50epds9SdHNCZXQJ31f9Hec1q3u16I9XoezpbT01Y11O/S
lFy4D3l6FZvb/JMaik2w0IgNOWUpUJRgP1YXfr1eJxAk1Bj5Uccu0dOXtg6phYV68kwWlEWPC4pt
8tQXaA4eLdDnz84wlMTld5KXRHMPwU/yXfS5b6SB4tYtAGYAKSKJxs0UIvKVOrk4Okh9z30Est5i
oc6p/Gv915cUU9NfxtHvFNVsnyIjJIQPKGKlpUKAIaNV0TwG9hmLdQFQKstHlAaxRxAk2pHycOpo
bH/vFUFBfYAux4mNGtxD2PcFz622CrtOQAcBi5QeRtAxJGE0RZ5YTtjjNhB7/6p1sjn6ozCKv0iM
RU5xM4NaF1VJbc7UBKQf95Yco7A+ms5FJqL4gaYj5T812serpH0uNpYSs814yJQWgWUgqUY5SBqe
FgibIirRPSj9dFuDmJqPmHvjxvWL/RcTtOQLzXiHLR+Epg7KgWXviboFqLRgqhNn8cAfkhIuGxXZ
8LxSM2nQRdB/Il8CMwY1JRvyd+Zo0wYqstjv0sNudcjC3vdZ3Lfcc0ulmWWDloSTFUBLd1Hu1QBm
7MKXBjGspB9/luE/h5eaYaLFdV86z/MFCn7xqMOSgyMV/7xKY9RhzTNCns0nwA6XXTtu5KCZyKgl
/0xSf2Hhi48KJwhAdAwNNg13uj6K+2iviblfBcjv2mrxi971Qy0QDYwA6TXvEtwSU+gHXsqeAR7G
qEDke2cU9M+FYQulNvSCusEF6Su06sibYEt2Q+QxVif02BQXN9yZkKfTIxKUlyz41rNFGxwMVwGE
U0HNhWWtV2X+MFe2nHnr8kzYiH8r/Hg6VvcvTzfS0iAMJ5zfH2/KaBNahY+oae9ivyasxrQwmmjy
nbqXsD8QWXN/sS/M4sZW6MNVelnggaExYdvOjQbODhF1gxX3eHGCk0RYZckpQvb874FDh0l29L3X
AdnBmR9VpsDjtQWZ8uMLzYItcniAF3hNcyRroyWOCPEul3UvlZ71mJp2gSB3TytTql2E1teB7eJa
+Ab1mwUdFB7TSrH5+WKWTbsnBv739h74V2/eZDJ+Aura4BcsJGMb6SxNPaJgMUqpGmO17+fpNv3/
zh/amUPV/zRye7IUJyYs5UAj89KVwgQO22RyheVJWhwhimIa77yRpcSIXlpoiUPMWHRo1jBCVVGJ
Pq5jGlf8R5DG3sbyCcwvgcbaIezVh5vFjeskc2rJ99ocEtiah/bkOppQfxQJhq6PobpNSVqIRTCP
y09nNPNs39IyA6Jy3sbKIsUvP7r56jGzOyTHd8RXh6+ONcWlmmTjKRuHvuLm9H6MTZZJAhixARo+
/8yhypocq+xZDF3JJtKmuOZd+IfNzsoVjSumYv4ZEKoMQvWK+wfgQ7gYpJ3dR0+nlgGBhMOFSqeS
1z5rWycDsB8rz+vV1GX5vU18pA7H0wqVJTwVsVLhH9cmWUnSlWhgvZ13r98srNCWVUFrIgxaMB0V
BSDFrgGK8QBHBNBr55FWuilUjt7fGx2QWCVpCMT0Jw08VNhJYw3eJ1bByYO6/YTlMffX96efl1wi
EsRv0/0TRlCid8zxqPn5x+q6ysIb2W7MKSiONx+M4hPANcLh8Say44ySQqoidp9wrbbmya5Pf+DN
uILFkXhrBrGvUf+vCB8wpMNVlAtLQWBl7bpLQE1IsiMB78xr/D5WYklzCvQNLExITspg+Jvc2d6E
Esrfx9D0VmDP92nzAuWQctWn/yvY8le8w3UcR2qRorylcKhsKYWjRO3qVdqP0qTtFxbbLZ723DMc
xMwKaM/ujQXkRd++zMxmrBQG+UdDd6e8MAtVfJjMSsc99pT9NEkJEhBCYJBUklV9uTSZ7J1vQRCz
OatUj7hye/ischVMIX4kPMoJsJEeQS47ldklOG9JR/Y7sLcleKkdC7M3165gg87SzpZvY5//Sii5
XhyT4+iMmDg9Ydx7XqhDD9e5hMWwbfCKMmMl19vNeTKCPDpESS8TyyJvBHjUbIaP4R+6Zt21pS41
ydj4VNSPl1KaB5meZXCJBe2ojKXSqWPx5TmdSluPgrM6HuQTCVPckGzwox+5GjWzrLoqL/Te9rpv
VKI6fZ9YhpXmkF/3EtqfCZpj3D0mqIk8tDhg9DdJpqp3/h1MXvb+yD0NZLAvEofxWBfLaXoMwrFd
3kiGd/kQL3BSqQTG1yokLM4O+MYZRgkRY4zSpE1vrjt5AJnWzvSDkuoi/NHfn6ujCxoAjJGhG51g
EwqoMOagMh64Rtg4ovtSGfeqFPsO3nyWUJXTlzj4s9YXoFpdbpmKsgTPUV/+mynJjaH4KquTi+5A
CTBtj+IBhRDj7ChmsuS9dMa50VrrU+TzwVBpjvjEiFxUYv20/+g5V8JGWQwmn49OuIVg1C+Y+svi
lwr27UG+YsP3UfVLWt3FeBLNf12XmAz58+3ld0LlOR7WqakfqnpnC3FASK5fdIxqWb7oXksZmcC+
Qh+XS2o/xW/hq4IhDXTUezt53BXkeAexiyMoUO5dwyiQpNZcxvwk5CIRS9HLbARY0cp3BIRmkEfr
GU1Od4cVUgM6Wh4p947kMAApxn6S8y++iApabAFgc45UvIkOluRUWA3G2jH+AH9kOYysN7fHDWq0
mOw1Q3mWazN3+3nNsK4EVozKq4UXnHgfoOIwW3lZaqEsPj/Z1NjenqssTa0l3FM78/ub4gRSf/D1
HJc4m91SlGo1KckqGP/UUy4nbmryAmNYOwI/d99I2/D972s8vouOd6URVoNuZMgx/6v1BZJcecL3
mA+9lv6sbq/hHh9iEprPP3HD6xrQyRImLeTcNIuRNDgzUL3znaedGELRu0xVdyiAnEUCxYHNQRUR
EochiLQuyQK7jBkM/se9OZ70yv86f3DFy+l0yDWU9/pywVasIN4U7aEGqqjFtA1AfC61lC61Rpdv
BweuBY2JkQ7O4mUkOuk8I5TKfkbl27hOdAfUGzSd5n45kMIVRfYxsK0UAP+GYOzBfTh2shH2bz/J
GfCQVBbmwLdxQ7w/IWVl91q2uDTmi5OZ1CUtc3+fvNKG9dstsaWokU4rc5kpXubsmDNlAXSP9x1e
hzMZJ6Z4VfgwIjiWmw0U77NguTzBGQXCx9X1KlXRoa3+U2QJPaprEneGN9A/LWN5CQ4aM/X8Ja+c
hGikkUxGEpj8FFIKJCQVYBsIk079RacoDPhtzC9FJT07MbCwX4Vre6QLrTn285+yWXbNTruI63g0
846xL492iPzfVLqoM0cAk8tomjjAcxwXXGXvFrtMAmSWEsJlHf/fvfMWneNvBfNJP9smY4yRoXZh
j2hZPYsko+n2d7A7opMSK3angTAIwCB0kosrydH3RZQSIPbwrriLgpjs338LQBzbGMRIypAej5Ff
lEmRw5JWCbuElvy20pFN/RraU6svcqBumbjKRmkKKpepK9qLh4xHtE8EYjyF5QUBXKwGcQOKHp3t
8BCN+56qZVqqQLrUBMcWK5ixApNt/Qqa/J8edUSD5x1Z+y2Cm6z6LLqWE/CedoJbOeZn15HSU+38
ZdKWNhk2upHXl8DUR18gV00HHo4/HkjMT5iXz966UMEYJx8e6GiuhZf9rlBHyPYswsqB20hVWnP5
gun0B6P5mQy4Or82bcGmC8fDFJ6i52b0iXpQpaNuSVa0Mvsel/dbwYlRhHbRTNiSLTT2qPv0TeLV
t5Rlwkgw0KPVZacx+o1SxCin0qhqhNUfF9o/NzLyZiS3ST7tTPSyUxqB7ib2VSBEVpXAd/llD2Ek
u0x/nKzDX6d1foD7goUkwUwzLixhx0AzyN3EDCMv1fEQ34BY3txk+3tfko1gcixlGbQkK0083hW5
mi/4vyAAiA/kh/6C7BjlDYTnYWRQbmsvlsDThwH38dNhWJwyqf/udA2fBd38d4xALFu+3SLbhrYm
SU+GxuCbLhLf68L55QtnVXvV9daX1+mXuds6ehmBh+bz0xsUj+p/R8B+T2AI3FQKsYg3j7hNOqVH
CHAFpaupKk69dLsRxf1h7KUIqGM+ny4iG+fxrWgKJU1s2ZpZ5+BMKwOBjk6b9VA19EovLLEHzPmc
PpWSqY1C1OZ7bqnpRC1oGZRUiwg+RkX0W402s1Rr3/VdpPJMWUH9zhUxOp37JyNKMfRCHayI82A3
u1gZrbiWG8ojfQowPUkgYABsbkiq2JskcequlRJYJj3wDZYhUD4qs51Sq2F5d6ArFdOGJk7kBNGv
IvovvjqkxzG+XYYX9/qAuL6xxbj13FWKWrkZ4tY4ipyPBLmyvwZcJ7TAp93IXHrc1SZnC4P2LRG0
/oVemtJ+1xS+4mcA3F0KqajaT5OwmZsD7QHeYpnBVGGFOcf1l41FJwprZ3/OaMEfuelULxo94wOu
OchQPuyqt//0sB8HtKIaitwUo+ghDqadQJTw8V/lPfJkObJOE55K/kbYl0LEEGUK17lP2M9rIxPX
/dozKBNsoA07pRrXvkmDQDy8qwnxAC3yxonTNOLNUS4FqKcc2hjuLMTRKbjU59n7++1ffbtG2Sqt
WgTjQhpDXkdhK03+6hN4sFu0Ue97y4tymF+31P4lZshLa39EWC4iwcOStNpdUYnkVoNv+foKVcAE
XmCURxBx0AAI0nLVoc47pl8GtZeLXinbJjmz4MskJeslYiYyIPPZYUjBobNiEbeCL6ZhgP4hObxu
kwv9pAf6kMylxqR2aC0I1pUdPLo0iBFbumCAWquQ8X5E+Bg6kLaQMMsFY+SYKIrV7p1NfkQb7NrX
RivnrikrgQnYGn2kBbIVVp6uKSCCjWzBJYcIseLxx2yUNr1+H/jfdVS0/8MKBvirnlOYF5cplnMw
zOyV30H+f9AskxzbTcBbKquxvIhJ0Kyv64rxtswiKpt3jg1mNwSbU5gT2fLiX7cl/YgrRE75XGzZ
L65+GfQeGCVGUg+e4HinKQOviwzGr13I5DQ7PyExWTZBp6bEc5T5bp/Sgi+ZPkXdM0McwfzPCOpW
KkOyLdzrWqkUc5xndQIWs7VktoVkr1vHNDkdtXLfYyLvfPBGUO0ShSYAYh/E/MwFoCBeQ0F98csO
QTRwIYF2KEcB/PcK8Lkb6lowF1BXxExNFxDkugUSjJ6Cdb6RF9wm8HQUgLz7a8sJ7uZpWZd08+BS
9JcMWOZkKJI01E1Qc3YYJvC7BknXe1n2BmxzNy7KNiFjKi/EbMWkeooLGJ+bZAKT4MV1diJZleOO
6Eioh/FxPQuXBInebvktvwyDn0pjxgb6wLv7CLraPNktdjcIQF0G+t3e/l8lV9yOSVuVIRXCfBT0
yWM5jHW0rdHVYio5iqdLHlGkc97L1DfgG75f4j8eeG2QthHHY5W2EWXLsshGhgJqj1R4/LGhBlqw
1Z1CxSnTbWFZMHvmakiqlFbx5NSDuEB0nQAczrEm/QwpMgTLphMFSiq6iKzHKYqD6Prncfh+KK2+
b2YO9lZxmezt68eNe6dX4EY5E7FNoacGCDC5qb1R+aHbzkYJRcivRtEaMSNXNcaUO4jECx7u9iY7
lAay+xEwZWHspT0sa8Slsqfxi9NO0+1dGbufTMNQk7e7DcwSXprwFwpFOC8Z3dwaaf/iU+E/nsKk
tD/4S61R6d+M7EPEO737BuwP/HbCNqKRK3mo8oGPU9bCO0Eau7ML2xHRc9W1kj5YxN1qtArEkKD8
M7RxHsoSwD+KAanybssG92GPpCZYJjouRfToGF/YgRW43SCevhAnZ5rB/y4RMddIj5Nncvm1mSwH
Gd4HQgfgKVA4yGYlmw/8ZEl1ukWy7hgY4k6EUK45bzh9YQa25KZvXB9YCw9A3J656FXmisUwVaOq
Kf62wCb+PydF7lhLlOVhkcmdkSkB+5D9Ihfl8uCGMLemP16KpF32ZeGCezriqCY644eFc5xKyClK
pxBoIHD58ofrSQFBQj87wrljiSm1qrbFGw0kplZej8GghHcbvq7LGlzakYhYVA769a2tOgvnIg9Q
Zf6iu0QpZMCHfAI2BoFVpI21wQdDv1r1gI4senlNbqIHn38zQAYSq8+SMsw3tIC1FaTjhEQ8cOY9
QLi4EONjH2kwITwvyP9jymeF81VZ8Q77ryvPIc3r/pff6e6O6xtKk0u2LrGJKiF7NmUySCGtJNAc
19F5LKm4qlapmZFxKS4zzu49jEyis775TY1kuRvSNm1cblz2haFMT38bAQ2Hg8guZ+EfdMo3BbRq
4It2LiMJxnilt9bFE8xNfJflQeyizlVQqZxrdhHlbTjmeQKNDV5bzqoLlw40EaFtSdYVYvmEs3qG
kwp89Q2dySa467OZiJcx6llnBjZ4frmWIxfMMLggPV/LnTR6jjgW7s6P75MsM7zNGv0BaN2MNiYU
R1ZycS+r+BLhw4ukmDuqfGAUvNVXr76OwTcaSIR8IK6wWOc6PnoYP477QQRSZ9iSYGqDj3+N8O1v
UEvDI8RCsJMOcwFkNe1DDnClMxyJSSvfd4/N2K3sO0K5Dc6sJmSjaJM3zqT/tlkvTc/kR+1hreIu
yBZ6USjsK9MqUKSWkuUeH1rHhVgeGipgkqcDcaiDtqkmp4gIOFzEfS2awZyUW8zFDPU8xwz/gGOu
I2Qm+aGEeEqU1Hv4PBxJXMNfcmOcP5nt0rbNxYSVlbQ+6zwskO0zEIGFTv2sJ21P2skjkYCnm/3B
GjSfY03uEAuGTRTxDzIOOKRtabuhr2TFrurRROLT97Z3MnGeeE+1HPXRJfu6rlfakMbjjtwUs7gL
I5bgPcp/q5Sn+UU8gvcitauy72EDHJ6JXgEGySKyGFFifujKsVpdRpkZ0dpwXfgOW+5GtgB1AdVZ
Vq0mxCbz4xp5whnXk1WKgEPITWm3herWIMYITdYpmmj6baphQ21ZmVJq9pVbih1Afg0NfTEkKnaS
HJLArYHZS0FRP5rtZxDEZXfQo5mr79BHP4fQkQstR9Z2Qzc6PQxRTxlzvQKTz23zHlAAPJpReE45
imuBBmTmhD9Xw83k+kcRWpQX+VJyXjE3tHq8cKHYi2oC0faRdMNjxfLwVtdg0yJPWM+JcQ3O5Em4
9hmSfv1hYhw7e1nYTv3z+S20T1R1bFYoo/vhcgy7jSy0wMBIGhiuVf7ABTKbvLmvJsCpHfPIhlQb
VefgEowC/3oY2eKgKUBnO5DbzK2oy6YO2N4kwXfS+XMLQEGsf6SAiumdMf0aKhZh0/ySSHonhZiO
MidcMMJASoKmznf37YL/89VZaglN1utqFckgnfp3W/KMfITB3EGYDwoGDEGdNVsSXsAzeGUPlI71
N3mxq/UyqIAmdLgfgtQgHsrnTWY2yjhq7AdGeYxGM93I8ka0iwvM7yp5EAv00vrFxRvg+n0idlbO
KvXQynOMXTJxHJJYXCfRsWrCwL00D72+Y9XbmutiSFbOBAr3LQqfZpyoLQgwt2OfNbLJB/KgkdR4
D5SX9XhnWgxQhEuzhGk2zSPU0Y6ZluPTZWAJGj4JVuIcSl272IePSkQ1xin1EVo+OJ5Tz2jjDZqo
JXhYaC0m6ygPo9dce03yBVmXRrrwg/qA9qzKav/GdHnh0ghkQfqXA2J6eppSu4C6WyjpoxDp8U7K
x8AXhyDZfc29obqgV4jotTiJb0ZMA3Y5iPXvmVSX+YZ254w5U3LU/79llM3sHxEYJi4ASR7BHHYT
VpY3XzJJ8Atpp7RSpA7EgWO6A3bUAq6cHMAN0BcnMntaC0EtHMJUfnuWf/9ICi9GRc1dhHYiQBxA
ISrdO1e4MbxQBMpb6mxDIz3XSvVS4Etv7K+/hNvO0LJCHcBd3c0za7f5l+KbHxFed4hFF4O6w0YK
9TCYDn/pprfuXs9iurcRtKJpN76lhfAAZMMapDKg9oHMv9066nFBRdahYPd5i9U+KTONdSA94kQI
zge9ICTvddhSPtHYYi0TAZtIqN6raxLKM2mr1giZLNNBkKvFyiySkgdl6qEzIrSXEMTLMaUD9EwP
ldyRLCFH6/rs8xYDaaS++85e76azUTXI9+qz7fsuWAYXmbOHz7KaDyV21tNKS4bs7jZvTVcaITst
ath6FAVAfmupngnkD+zW5oFMsC4VI087Q5x0N4UWDuKvn5SD9DLSlr+hVX4AE4WnRCw3ahqO0HoS
d+IuyT6/WQv1sYcWeJPbUVPPTIrKIHl0pOaGK6IoOgDYhIfoZwLEYgr45g+xv9iBoz6J6V4zDzxv
ZY9oRsx9jRz8XE2+7w+Z/ZztJOkvL6Em16uloFBejbd7ojkcqr9WqMfdy2tj/+0pBg393Z5bROot
aseGWRhJ2iMWhVgLFZS7rh8aBDCGKzcGNInefq0cLRNoSwiy7tBFN+XrOvv+AS26OxUYEqYdPry+
Sq4d46jnbDTjQp9KtjshdwvRirBLBgwAm1Rjakj7ccmIa3XZOW7AFIlsf+SYrr/Ld6nH0NEA8AkI
DkKXKbyO8OkC5+ugw2G7kpSEL+u5k6aZgoYotPRjPilQtJqbV55rPBsAoTAg9dtW148It7rC4SoE
Fc7OFvPtPNvcs7+8DJpCujAHKIa2mb0a4I7K78ayYl0ho2UQqCG4AQQe+hTFcoL+1AblFXFvDEwA
HxAY6MJ7QvpYNkoDT0TOX6ndWkcVrisXdMD438xrh8EFDphQ4cgOflgTX0foH510vjXhMLtRaYuQ
J+y4Tvf5qYtuZoDFWGrMywz9VMEn/vRShNVdIUxoh+82tfBA2Hm8ckxUTHiTu73RlPD8ePHV8tLt
JqYAkJy30/BNdL7yiRBWGTL43V28q6EAVMeWCoXhD5JF8OIX/m/a5Bv80hvmuxYbThbbgfEuqKPQ
9mhwV6klXZ2hLII1yYGeuyP4o1Pqj5WU6lOTeW3Xd/6JLr2gvn2Ggn6PONTQ4M9dUjICSFWAHFev
3qdg/Km4EVpiNLNnsfq3AMYsIfQgFv6R/3LR3XGS4QzFdw2UbpPtBZO8OfMPDvgweanNH3FuIGSv
0mfq3SI59EJxhNxHz8VnBWtqH6x6xkJC9ag+rXfqlUH/Mpi2PqASnl6JKoRImOYwtqZ45r7SwlPa
SwHb4/Vz1t387coSnhzDWfgwU5KsArZaOXEF2CNb+jQz0iVhs2U68MQwF6Usja00VR74V0AaBP4v
80aPo6I/vlwVB+NnaxnX2SbQIDeGvy6FLyYhiwdgUtFtfIz6j/NQAB1x8cv1tiSE6Qxtc6MUNZ6t
i5I4e7X2WeSAR6bmxhCNGFspFoBvxJNi8UBNBk/GG+ZJpiIdSoRIzOJsBFFIfCkO5NS32oNc1/IS
0ohvESirPrxVgprNsIjK/Nf377efdUHWJeKeLOHeHryTwvbXtR+xuQTes0NoOYuXLm+UxTNAM1W5
qtV7sqKZmvUWsb9zrvD5MOgB4xiX43WJfEk4WZ9jAppKuccZ7uAqZcjB/m4pa1FimQP2c7A3TDFI
zxQBlEPV3kR0bdcL1pBxIofkeWsIKYKVNL2QKsDs00+/cKhfbpu45+msBryW16hoaTXIhMIikWs5
m9bN5hDds2sthBag+4dS6Xh/2Baqf3gt7q8sNVwgNUoKcHAEii7OHHCjlEoairZcoH5aZvxWuBAq
FqK1nBwfYRvLpblmBYCZC7rtbr2anhCu7AZRfACQIvb+ftLwemSA/219GngdbbfTieegZpiOh8ny
G/OSLlaqihlGmTz+p/W6VUfhaiuULM8FjZDSmLcak4WLV0gE9//sD1pPPii3CGks++hii/Lib6yC
snVigY2GTPwWwjro3EfmCNTp9wAoDePNCHOQdsG1A8yN6ZEOaXlq5w8n02hQ3gbEY8ljkuCj9ISz
p/s9fa7LLhYKbp5xBUSKe1w9zbKbrwxKfQ6Xq26aJ1IIf2a0AYv1zumWP2aIM20Tw4g3fDXbvMQJ
tUd0J2NwE6rJUSxJu6CwJeGnIkUmriAf5oRk5VLhcySAXIdtVc7dmGKfxSebLSM2nC0JOTG5RE8P
DfGPoB/sZqEvpEUZiGjdmcVGxnsSMMp9VbotnT5GEuusQDvgDB7KfJiMd11x1w4SAuQE/eNTe0rF
vP18B3REhq2V5YP94u2AiOw5CcCOqYQlqqriuwv+vgLIxEdHnSz6HpD62H+ifzkUY2mhH2piwAwf
VOVhsyY7q23VkcvQgoOelw4ZhUoogYQXTy8hgElZgbA5t+egIofgNjFCLHG9oU5iMCiETA1eb+OR
s1SCRgcsgIRsNRkKKb5miICvnEumkiHX+zRgKq4uDQRB82kJYNc2wCRKpwwgSIr15Naszr59cmzd
RWfYGRmcErZPrUE9/EtpqvMNyfPQT3VSBwEf+yPLg8PfsxTCOO0FL3BISRBqFidvUT/tr9G6WNDH
rKPsS+Guhq2RJ1+4Jf40bLQKaAdn7ANVmZk/lWGroJpubsxMQ5ORFdhItSjsvwwm7WTkneqL5ifw
eOCmbaua1oYnFWt38DEJ02MHJDihHBBhwcWuIQoDsMqoMssH68IVTdQY+s42Tdl9baFfb868W7Tx
bTD5Oa9Rod/7hY0yAcu6FURC95I0yy8d1LLeMv7Qw7337jULHvG2i/w5ESwBkBkdoFkF6rdvRjbl
oEYqwtED3skPs8GdEHnfhJ4nkrJI1DtCp2ZOpIP2aGTIBa+7ScdihyZlryBrHdL0RsCIiP5rS4hl
fKNcIzf8X6qleB0jqIccU085Tj9htvGSkZyLq6mA3iSzQn40QyIua2+mPWZjygV4pLxw8IvvbnjH
wZvezKFXKMAab8rRITbgYMqGegQ4l1RCIoHzU/SVbN+5xzvYl73cVSKWEYSJzCOi55P+kc+fMHK+
MDUzmsavzr8EEsZA6F+xqKidGlwWD/ZptEJTIVMLejE47OmJWxwfV5jcAouxc82IZDomlg4mpRIi
LmKN9ftCt1EP5QhvY/99rL4NYq6669jO1qVfQaG73OHSUVvOEDCaXqsU6ie2h5+Y9rjQTUAvm6+U
XDsQOHQolAw8uvtnbY70jXpZPtPtcXAZTqNIDVhV00vAVATvB2JXl+U4ckjdtL7vCDAGZg4Y0WGe
/QfSng2mhnTLHoAWNMPwpVwxx/vHFet5iKbzdhXnsM8Fbv495wU0oQvj8nheCzC4HE+dzzD1rCVQ
6T01r0xIxM3Vv9WzEo/IZZum3+4WZdj3k1j6bblSsiwmyGZd2wAWfeFXNbYQlDhx0YepfFzKCyZ0
Fbhy+NMw7//7hXaAYLQMoxomeDcTpEUkFTjBtVjZoLWcM9k+LgB3hv9jTlfjBmB5kM/X+6Mh3zym
Yk/3sjqQ284Y52LgdkZHrBsBi4ehKvCf8p5LJfzawhxX7NTjiG4Ez53xXr0pp7TgYPv8LARv5IKv
Ftx2Ou2bBH4CMQUheYAXPUZ/n1v5LkrwrWs4nLaPunWzAYzHpTZxRNDsMNfvFHofuk4zWTj4q9rc
W1TaWC7RTTtU2IWJTK1a2adpXGas7AahJpZCJyQbH3zw3gvTTEiifmSIk9UgFZ1sHC5su4Th+Hji
FiWZUbN4OMfQS8QnMYr6FZf/yZ2UdLEHTvX7FN5dRvDVD75iSpWJ+HgTLt8DaPi9Qqj/W2FuthWU
Ik0uYTz8wSnG396/BV7sekrO8HpdR3D96nDq1rYm5WD01uAgc6kRbCNWu8Rhp4/XGrAb8IV3RtSJ
YDaRgBsUi9elbIzoJURo8suk5lvyJH7S8mIXPJ6ZdduNA/IWfKwFtxKSbHFd/W+wL1mROTrNo+Jo
XIbVl9SJ8sCadRHo+AAHUid2VZJM9C5o0g4y2s6NT+Emd+6hU2/4UeSpoKpwa27Q/vw0GYakyfCZ
vVrTFzEwFtBvGLdeV/g67tEWGuskbDlIfZ8oyGaCSmsDXgNjOzP2ekh13QzlS17BfASIuheaZBEh
pw6Q4fYOvwsp39giKg6pQkM3T9EDzr7gXkDJOzK5NqPLRmDuiV0Z5We8DvoV2ne5WI3HriwXSEYL
2dVu+lL1+HBjR9D7nUYckjbNbj/Ra2MlwltXqtu+m9bFbmvzhLdG3neSwQWonFBHjCNiNIp/J+jB
Iq4FIdf4ACidUyb5rWPoqIaoDVuRiXPeyFn1oqKT/M3LSk+CQSrXcYSbuH0ODLUKTH8BUKwsXTrz
JdhR7n8cG806wep5ML35SCDwDxMwIutbXtYD02XSrM94M7ai13m5KBD9Ts7dmkNQ4+0jOERJ6u5v
RmbfVFa9H8waLOQoZxvP1unQ9yWGQU0Sc9smGjJFzFRkb4+BxeIY+I4Hb00FWKN/LCHudO09h5Vf
iwQ2bS5ZjuaeVlzUjVxQ62axiUPxCGLU4E0thQx0v31av8uunYQHmfPYi3BdYDn9wd142hHshPtl
sbes4pZenRePKJ3DEUGSHFNs8RCFWxIqMac5z6p+wJl3DJ4pHcb1WeDi7TJJiO7hpuCvuBA9i/KA
VikblC13Z6KdCHEOWsKVo29+jsITO9owG9p+8wvNqv2FdpUyWCNfD9iqYZ6bJUti89W5FT+HMZwQ
jZ5mxrHcu6bhWf4DDl0A780qyTTJAL0J/VrtBlWhaTeih4GuHP1jBrG1ll7N1NPeCXNr8WAxdSqN
Z00vHvNg4dw61klM0VhZkRPSBobHpt/UgyVlgJGKP2tO8Hx97fkQrS4Nv7evBcsPoqiz5csnVaLC
l4av2yt2891FkZB8CNaKQiBy02EmCn6pzY1TZ2hbAwpvluLjtbZOgdPFZ0ezmm8XeP60eGmVLftF
UeB/xxQfdrVBygYT0pThQbEamlH5w6OUIRPAOQNqgi7OzeaQrdQwemMwSrgLbcEjw+mDqzaCZmpr
j2odt9YbR1HKktLTrV41UPCbGtakzoKMIa/ah69XfVBHkaVXYjjZcdQAsuH+/GwKfQB6VocUNl5/
akQsaY0TfTXCnAHrIm+25L4amfNiyB3mDieivC8MSJInLfOFd9zPfVyDIO+ZtknBNxNFeC/4/Oml
f3Q7luL9RQPkyrgCWNOY1Ypb0MYIHXG4IgEE+BB+zKLo4x/j+FFi91m0juNm4gUOKpiHXY20dAs8
rjO1Vp9KnKD1JUaH3AWOSb5gAy1R4+1rB0uC+CRSoCe0OPqKlbygPiMdAlJ+RBmNsAoJmbl+O3Ux
uST6mv5hDOAEuC72sWG/uF+l6pMkTJT8ybneUJiQKd+tPoFVdtlWpCNQO00J2giHfT58/wwUvEZd
iSsouMnKGbbbZXEfMbg7780QfmYGODOG+iJcZEdod0F3FEh6GpsN4zOFnEmCDDKeRfadGa3QJD6U
r8DSUIPYyunIOeEqDYFqRt32bdSj8vsi2JHki9EJet+mKRMqpWCleFutov8p2Fo/kus+7OqDujp/
3WMAtiDBorl2Iq4bX1WZbT3z/r55L2RCy6f5S1iTg+rwYopvSbHh2e6KV16VbLZxpCfvUVCWVwBZ
K7I+bOsGOormWjzJMzkq3NDNY+PBpnP2COs4WPS8FTgpgzgg9GC75jVxXyP+qHtnYFsxsQu8uy3T
dOvUN5f8S7khIAsWcVUFM2b2KF+W/MPebCdOXhq0yhjTlRu3FhMa0JqJh+7qN83r5k8jy5ipsv2X
8oqXcptBrqXQkeQ6egV95r8gC4UftkEFWXK2U/4s/KphOc3IbcUZkgHMbjCsPPcu6DP8J2MdzDoC
LW033UKZRsVOpqtGurg+qp/WD1vHzRUubT53WVtpjjdFokEEo19OE4uWtBDY7pIKH+TO23jjj2l6
O1OtD2SVFT0EN3ukIbalFDM6/Kwi0BzaPx3Ll//3vFEX2aLRxFMvQc5lZCk7uF6B2mXTfFCARzIV
ZCY1Y4g9SxeJICKtm7+AtRF8knVpg8v4jC08pECmbIPnYrwin4TS2fYXJzpdCnSz2Bz6xvJgsC4P
yQryDA4ucH34CC/iVgPo9dAEmw0/2BqXyK11+7nLlXsciIQP5cO6Tu+1PKh38tTEi+ubIqgwnNww
rGqw7VPDwqSVnyOVokHjE4+hGNZ+xbbPq6myj6xPttyKGaC4P2bN7o+NU+nM2VyjWVW6/ObC/kjC
wkITLI7jIYN8FIYVVgzk1el317TKCm38VZFGCRD1uB/6LybKDfyqKNVqomeTaPr4AxnA6vk8j+A8
tygVZGIAafHfuTCS3BJh1WAR1n08kK9VocEj+mWJp/5RtzrSUbEPEpQ1sbZMaRLJPgG1vvTELKE8
IHhMCmDQZm/RGpLg/rBKdk2MM2yOVwZVfI3I/oc8H/nLxa4u2oUO1aueN+L1CWS6NIGH5Byu+S7Q
63erCwhUW/lbOjn1odab/0NV+LOc38v4iSet1e7guOvtEHxSa+sqX6dvpWbBINU7XeXNHZnPe3cI
SmEs5zlqx1cfnT/JIreQ2qZAl2vjGLBcgB/66ZBNiWhaZCvk3UNbY54Gq1CLFSzowwG0TO7MiQjW
RCLszM29kRSAC1dNuU20jYvmyMXHkoVvHulGeeqbIaKTZmn3HwEXCHt4y+C/xH+Fagdkg9JJuyJQ
AvbnTzVDiJJlVXKknYFpqnaAFvv/3tDKmTwu6i94lwwlVlMtqa95/7b4yWI3NhbDrh27FUNA1FyW
Y1gh15G0BZ3l5xrSsK88ScyahRuyktFrsLj+FcMbVlIIM3mf/PxLbH7qk0EnW1Yh6vc+rRiuUACw
1T7H29Sjp5L2uEPXpsV15cNNNH4FLcKqrdTZxHwf+28epIZJcQkeIXf+Nrj2nR9m32OwCcp8ZUtt
pl9Gj1NWoLh2oGsOhpdLnI4eqbjIgfTBO+MPsfZTkPwl/8qC92P95SAz4VfWjl47xaZEROrITchB
a4yC6BNku+R9x4r/8hFErE9zjEaXkiaMg1HSo0m7XKySHSWHx0rB6HUNGmCfszBE+6eEHpPmMA9P
8Igt1i7u0n5/BTQGOrjvl3QJhzZpxnVzjnpObKyE+A2uYTgmvjBpnaeWpd8LUDxjUP4gctDjNGcG
h8LRNT0n4F7HXTzy6mOFt/cyxTwNgZY375nGuTbFZAO6RtCOXq2KchNabKN4BikT8Tkexaxf7+IZ
e7Ya0g2MJ6DI9wAHGwmjWH8efpDEpHOpVfDBxDAo1cLdRCdh9S/N3Tliy9IziGPSNIzhXTuI5ZV3
5xcvH8IvTVjQwabgpIg0NGb6h+5LtHRpFZ937aVEJ6Z76iI3pMoci7LY2c6770YrVTF4K7j4x1DX
IOw/a+fvoGEIGyh1lCAQLqlT4O7RFBO6qD33qMkOjd4p7SB3Iia0JPOszMWEbbCnVZRDn27nUj/m
YRY3uggXDPONIaLDnA/FzMcLwxd4UGi40mLb1nL57MfloEuaLvK9uOmRyJM/MX2BakB0MvYTnYkU
MrNThkrrQReXWdUqc+75ewwDH/nA5P4dvWk0x1LVgDpMBcI5Qs3CdYNLOhsKTJQ8tY1dkMG7QtLS
1fx5SaJC0xmyItQgYF6rZ5iSaiT46UOBAYGryppCGuQXUjGBxLt12lXKOeT5fI9vTTk+4pvCJOau
YyJdTzb5Xj9enMO7DkGjafnOVBNmTrtAoVrwL/IwxAKGIMhjal3Z8ji2Y6WPKqr+9IgNZZTeiJWY
sjw0+efVITfTZuEkHjhJ4wDydFVQ+xPLrgFf90AZXv5Oc2nBt/WsdHqiJwZvG6FwcHSOyqAUBT1I
SPA+UwIQ5+F7pJjOKXme2JrFt34r6VlPRiWW4410+Gif1AiGLQ5oWryD7aV8Y2uHl9V/vi7ivHxD
ME02ZEQjmrUMJn+3deCvS8ebnTVpEVoceKcy0CxapKKE8MIKpEeU+wA2IlOHcLFp5+8OMJYuV2Dk
g3M4qHhSlW+2fOknsXJibLEgldpkoSvnHQgB3trTaYn1toFTaSH5FHmAdtsWeEWd3YtIwvednp2d
3lMYnkEA1knocCWzhl3xl3k+VAUK1xXiRgMV7t32E7DOPt/PmgGq7F1lnn6rbnlnkMDgDZC6XQXB
gecU59anNzbh1TDIO9YEXh4WIBrTZgTufssjaBTn2dSM9UgL0bP+d2bCu7FSQkV5iF25Ccq3nEv6
aMYaE0uT5gSDjqH9YjaS8zAaJCchDiGJt1e8vDNByYiG/XugDN2h/kfZz3R56Qye6dNWMaSA4Vjl
SF75s8d8g77fPad2i24uirS7OeuNw8rIaIm4tJdfXr7Raj+HbflMztpLxQUsRG52wgGLC0y5vk0g
Jamr8fKziGBGNMNgylaz3ON4sKfxyVcH41dgGebqgte4zsQBPtZSNdsgIP82z+kzNlSqPRuUcL3u
WbhNAhcMQJvDrakIauQhTorosaWXFrrdzdKVo3VwIv0mZ2CFEsYFk9fDUlaJMIKCyO2taDU1rofH
X9qxwbZDZiTi87ImWrYNtZlyzViG/Zp1CRvjZHvFJnKbU7IuhesiV04pNrmI6Dk3MT+uOQI/pmxc
uqHs/A28JPb/DxyW5QlHsChnrCmEulzdOgAFGAXq7aq5khUXGWBqtFlikZ5VZ7IQLRxWeak3RPHF
bZ9fWcMAPHVbdtdWrEu00Vpd3rXeOABST42CLPTZ1mTJFyPcwxvzTPzckCPi+JvxNlGRBbtLmArN
ucZhOSYnlyf6TZZ7wwLeux6e+BEaVYln7ZBgN9gDa3onOSzZ7x7p1LPa1vv2SBk/4l9MEDH0w/Ne
M8mKnydYoqyE8u1iQphGZSrsC4rzRJtNxQCvKHqnPStThwi+0pA5YkAPx2tL/Zqad6QD99PxZRfT
Rg8cgx8NiyyGf0sfZ90K0rbhEfQGHteoiM4HaRyxfLr7Br9lqGWeW08/tmM4FerNLRQ5SiyZc4Pt
MwWjXf8WhXAJb0kZUfVuzo3T1gUCNqCTyhciSYxGaWl9rbDE3PdPyk/UKlfeYrCgIOD/gwKOHfPj
hBmFk9mKlILH5WHdolzqdFrRUmb/KTTlo0pQ1pRofzquXzOUzDP663/PkC9JXUWzJ/hOi0twKHzL
kFxMEgfIWT+Dcycd+gzqCMCN5cERGV0+n319A/V3MlgAc1ejOf4xSjH+WPGB+OqJZduvKIbhgFCo
+niFZ6rP5J1YRxhMQK63R5khtcCXUnnBcvNBducPxBHNn3hbufu6nTqm4Q/K65DCgcLeUQK2jCfM
jhm7q0VQOhkomKxgRA5QzXDQIXTHofNDBaZkB6IUOeBSFagQhcvZUpVJg/yqFvSJx/fxe6g1bg+5
F/AwPVQPxjnT+6nrgeBAxPupqf94x54o3QyzNSXKG+AdaALhHQaGQ+UBkIB1+cqxNbR7UPiw9lfc
cY/GWtapThJtTtBGM02bDbnB/eemXDx5u/X52vvxgMbBMuQi8m/zTSEnTln78BCY/SFA5acth+3O
kLZ29rCQubkbWzQmwN+445WLbWGD6VbjunA2opCn5bTKqun2Xr4jRSgls8SqomNcrC+SPQq7frwm
+6gblgNCSRLhGB4mGrYC9xEf2o+CLR8zcAQkbde0y1FpievuggSLWpzBWdW7xJSU9AEF63jItjta
E1Q/PWCOefbpYd2+4JmxJpG3LTtq9lYeSsPcofPLkQU8v38Mg/CfuVyNj3sSdok2i1MtV1FsuAM3
aDXngIyepvDlQ8iebyzWEHzbUqWjKLBkOovL4wxFnmstNVFqdzlCm7LGKUkDQhDLovuidvcR3VsJ
byOU4Bu+rpkbXcSZY7LcT0uU0o9CXT3EHmdy+dX1f9VB39xxxRutFKFctNq7+F2axn9M/m+1HxOe
O29W4a9JVgPdgb4cjU3g103OcRx/BYFqsdVU5vXWHkosVG+mrDZLbVCQgvs3/KCUZ3LsaNakdi6Q
E3V7ALyCc3JCTxXsfAM5vo4EG8gQGu5ySY69HDUj44dF3YY3t5gdptCFIvlCIQkLT5+CiW9y/JeO
DEW5inchveNZz/gG6T3iQoj69b9LqJUqWSftHMAqJdWSAD0laRlaMBmCyKj9OMuUKHNhU7xUWzFo
q3J6zu41XYlu8AobEl48UtDoH1GlpJt+MXwK579cH7eRM243FlZvj691U60SoFj2o3tVDX26VO4g
yj042G+9ZPuTAOf4F8lPjKRpI8lU1DAIkbaGmG0JkGO9+fV7v/tDgF9dOBwpP9PT/p5D+PTZMB8s
OrAtHclVrgltaj7lOEGROol4RxeCCndi5vEvNKSbCCTQGoFftZwK4PCzMKUwz+ApMgC0alOEF5zX
OYJL7mvs2uxIYxlQS+4L44wBIeSxAhEXkehbEXHOJsvlnbOkn75fRKaqYYElt0s7CZCljcheYhUr
GsNH5coum+ttkHZ1hvCx8IlUfE90KCoeI49BQAGIMbqK2HW38FUKgf3PkfohpZ4+cICdEKuPP5Qd
XISYiSLmn7ksTgJdIAE5Uykx3QtmFpqRVWC66kxEMYB00sXNlK0hVQ1w+VVQ9+cKofdAFE0Jjqk+
3QRrd6tWuEe3kRPEGzVktppxSaGPtFU8+H6xSwW7ZjPPztJRcKmVgjqUjrC4dV7op8imP0Ne61i0
9xkenHzK6eMQ7TTw8GHetE7bGRX52HZu7BPo80AjWvZgON6zfZ7jD5YFQMeizRNJ00vKexZ+nN8S
huO1kig8V1nssb372jymNwnWA2k60W7eN0EFjvZDYmAcoeg7mioxjzpWn0j0siGLUQXrGipaWqJR
UEUpY0FLwLSjrJEf2/bHa0Cjei2Zo+iBZrp/9qYo1qX1HDhZHoOzYYBwn38StQcz286xpNK1un3c
4fgvDleVpAJ+KpkvjpjRRTC8FtneQEyHRWA1ycI1MukfEqu+Ewd0WIf/hmb5cR3naU1PZaMg/B/X
aNn9DI1GlUq/swPsTniFNeiYIFzmGJwGUhFspGYe7puS4meKyqCQrZAD/Q3+tfK0GONXyH4b5BEH
QuVt6WYSY68VEo4oGmI94pUepjg1Y7kYzzqGycPQaMFDxZz9Hra89UxVIP2eodO5uW1z02vnK08T
wskJj6NG2Ry6BuSshPxKDhZWl+Ko14n1tzRIxZRnadnif+W28OqbiGZ41Ndg0/Xv3pQUXIeB6SdG
9STzze9hxLW/Z1V604xR/35j3/MYYrzigPMlVs+hVcGpp8nMQj7dcULrFkwkZQYwGwr9i9gbFUfF
lTaaRwJpl0CulQ7RUrD0YYAkzD9o4VEGFDFz/2GJSMLCPoDYLGh2x19R0VnTMttZYZXTyh6OfzFK
yA3Z6aRIlU1Wr8w3W/e3HVo8EREVnzVrO41riKtfmZiOvUO7rz1umxCmxgut32qtbw60rkj0If1u
F2QxB444/FomnvN7ACX7G0W2f6ICziuW4plxOIOgWybY37EPDwTZG+PvPCWXvMtlLqrAYD0P5UCl
a+xmyDazcTictVCcM0ZxZ7k5GH0BBoLP2Y/dSBGQkVkL2H7Cmbypwo+XXuLEkOxQYjr6Ss6wZgke
6j22CSA1Oy+2jFd9hW31ysjGkpWkH1keROMmSLpZAKLbEYybTPkGzQPt1yhM++sBP4jUqbLyKMUY
ji8iFcZacJs+JNcOM0YqUFO9gtqqTMmVJjzx4fIwA487QNXGQyKRIXMw2/ksRpoxfFPOe5a3DUTN
HG+wfISb3Sxm4AiJaSIpL34cldjMHiLgEZ26zQPGw3SAMMrS4S3T8LtSODuYSIp0DYEd+u7LQDas
1RFfbp/RKJ/fQHE0rvupmEKK35EpG5JxRqSvUnmUi4u1A5+9wULi5iDqyxma4WYQ0/yIKL1ddasR
fpXTB6ijHrE1zvb8a7o++efA386LsRY24WZw0rl+DkO2WQXXl1CVaf99BigXU1311db4KieGqfbT
KUKcdfUwbsACDckB/BweITQGRyAD3fQKUcaZTFALXhRccPH2HScmWNM5/E14tZQExp23mT74GOCO
t+XKrevHpzwaSTx1XnKhtRsE7OZSLOXErmYPCNXseFmq6IqlDVpoiE5cVjmZRa3xkrARW8pkkSw7
TJ4DgFjWWse6wAbdVelYeZXu6kXtXuHW6/vVdSgMUbkpDqgxVjCh43b6ibfeUqKKaJXHkuocdC6b
g6g9G9q+nnB8TCp5XXSh1oGWIZV0GtJSD61A1CckPoKTbkD3VatLEQBD//C/B+TCWNgjZt3dzXsB
6jv04u/27L1vHc5jHw87GXTPRA7hvZwAEUNA9gQds9muU7fCUSN9z7q92K8XxqtC8g+wGEf60Mns
KShxpZYgNmyzlnP9YCmRS6J8bQ62OdJLhucV7Ge6aOpUNaEblaDtkJoLtCmJdQav4sCSZkmeIbYN
iMEnqf4RhjPOqPZyRdmTyPAmex2Yt/mfloyGUcH2nfCpj/BxA4J9ZBUjC0pT01/txrbzbt+aKewC
YFcK24Zv0zgbOmcwC39GgbI+Vsutc5byX7zf0VSP5psihkZ2MyI7Xv/zKwQ6x5wZJN94r+X5NKec
ev4COhec5+KTTQ5ThDRE8nHHnFo+2+3GXfXyEnkYWdOKxESsUt6UpVwIKZjFklNw2Quu8WH2X76P
sc6tffUGTL4WDWoaguJFNDz8N7DTI1TV0dxQdQGhUhPhtaeTk0/oeXgQWorg4pSMn9P/nOvyOKzF
ecY55vQrXceucv4d7gKbcQu5GP1YJHZgFF0zTK7GLW01iTemZCdAvUGNsHIlF81vyOolPuRFOEcJ
UINa90qpPQ65yVW+mrU//jfj0SHZnvIVLxQjJpwVaa6TDo+2N92Ud3206MxM6StLWTCMFRbiNrM8
2YQQOEBzUiFbzn0emRTS8yMQ0fo3kzRWHWuo8UFCuT51sVCIsW7oQ96aqtKlyphb5EDLDyQxxqT3
CKjaFnvdOFEH5QleluQLZwrQKa1Tz4Yhr5MK1wBUgRZd6akxeRTrq7e4TugBfB6T5DgUEqLo1Nu3
dl7NTRn3QWhjI4xBhOWBJz+0iUmBkEJaRUhUR8lCL7/r/H4de9QFQRgO34bVS6exjc1k4aspZ+FC
OtE4s3hcziwVnWyu5QtCA5WB50Q96h39Q21ygXrEZ7pGChvBWeWUodxR30b89hotK5wksnApFSgr
TjvK369i3t6v1Z5uGyJIW8wiv/e8U2T0pzof4BL66lTXzK4p5se2YcInsBYJhJ0ybF6bsOkoxHpr
bFEV2JyLke6BWL+0gsEuBW+HwJaRML9ZcavJYpB1JY1Z+ozraIhYw26vcTnsaUcyMaHG1v2/ekWd
xlONmbPQjndWfnzQhwT7A0cPAA3uOhzn8qmhVzAXCf1IQMqeQB4Qe93sdRNfijBphLMCBW5nw+Yc
owN8XFXhPzeOQPvY6weL+qzLnEOW71FUWI9Qv0mbEE6FV5rk7PoXRsq6emcTgF7usF92/AOtOgz9
YA4Lwvhu8owdPPHvMA1r+rhMuG82TB3A9H00XWxE55pHiQk+uHTq5ZsluxZZcAJiMYG4ZpMtyO6R
pVH/XsnYgtqThiLnHlBd0XUc6d5DY/JjwOstiNN3kypA2/p8HGPuQ/SZ0mJ+cQ70USPNES5QeFUe
PhnIkzswaTSiBbobsGcDIZo0qigw4cgYMlt3B0kdC4uuoHZk9eeGujTHgE++Oxl+jasSZvF91fr2
F+6HKlXzFf7p+9Sd3aWF0NEJsBIps3w094eC9ogX/6vNHDjmOZKEHs/qAeDmgIYkpFLvi3AvqXTl
E6dvEba8iKW+TK7uocuhAIoWabxf4KQmWXg7AYA4keWxhDY1r4wPK7a4I5un1vnyZB6TyL414hIV
lejz7ag59H11sMMYdaT+J2tWYyp2AjIZ1yfbJ1n877PMWkIsnrc46YmAdvPuwQQINh0Wo2uHgHSY
xQYYxa9gA4w+toquwHhwtHE0mjCJMKbz+8MdpH44KdhWNYJzY0RGRbmNyD4ucCgIzVXjK/SkpmCI
xRi5wAxwI011K1KSGzuNJmNIox2S3SmJmNSl0qjVb3uNiZIHTkDwG1Dp1DgjVP5jiqc4YuLqjDj4
iGMRMQfSPlNUHTrm5Yx8bkVod2qGl1zlXjwVXNRJqkaGbYG19qou944nHszBKP8zW/BtwyQaJFrz
6oYvlwseq2Faxs7lGpDBMYsGwS9zdC7cLxsF1psNIVXFNcv7pzQYoaGhftav4qubDspTPerLT9oi
O9o7oxNm3LzkuPQgYpvKSgYupqRiimo08lnHHpsNiiyG0Vo5G9v3o6voBdVn725wjAJ+axaG2A2Z
9dQZvNmJHsz1W+rX8OffB3l4Olk5OeCJ5eT4icuaQ1dG5bwJE+liafjb999YMoK4Mra8fE6vPYUh
QlwazbUqImHW61VqRzKyQjmqj0dsm7vsPC8Z3KI/Qs5rh1REt2BYlQzLJg12+GOr90vYZZaN/TP0
rFcheLQ6PxpFQ2bARA+MQRTfJpTTcHFBR4TDIVB37c1F0ID9qA9BMTJspD38BmkopCiP5EaEY1Gv
oe/P1DIslrF8vUFiwJ5W2kzS+iCZsU1FXUK18CCgE/zHt+X0c1ZPWIbmbTPPKhX9gOyKs/iCJs7n
C8hKvaxy3G2xi/MPDAdNamzGUq4+F6oo5I6rS91DjZA0mVbd1tuHMNtPx5xTVc8B0VyQcCUm0Qid
ZQhlhprQv3Tpwh4d/Zx0qgijtcwNRedFwwSx+HmB9yYD2m6srMAJslId/1mFellDiRMBVlRdl2Yq
xOjCc4xV8FqdXJbpDL0HOJfI702wSY/UyHQVY2W2iSNa1Q6ysUhNkVpW5az7JGnXnq0Ep5+zYGjw
FfT8zqi1GFKBZYyI/JP0aU4fRdfHt1nw/7IlnaFaVLavcOcEgR/PeRryTgurZvwPktL04ccdxjmO
q3DAdedWARsLVEi796DBhTiQcexcNcV0jt0k1Vb/tEBCKoG6hH+XxPQzdkUjnYTDad56QeaoiOvW
+25fvJEtQZsmTESn4qwBeXxbjt7EEVK9RuFTKjkRclJ/eTClrvx3qAWuABzG1I1Mz3UZvnBbHJc0
sn8FwXQTUs2P0HYSkXVhaX6KDhfaSip0nugXAhbbYM0prcjMSi2aMc0W60BAjhqNxdox81sbRpM1
166Mj+uAOHhiZ3xwNfkrGcTwnatKqaFPd9oIF5RO2dnsnQXdBbNpXe+JKGcC4wZJW3CDp5MOqOYK
RoPj6gLBEtuh3jthAEfddyckuHhpXWMr2vxlhXZezhX5YPG3R+eRxMGtmRruJnVtJ0N12p1beVux
xF0vqjjS/wyRQQu/eMhE5bRox2mT1gZucTYfEQLidIwlGTA26DEJPMSdpNgfXJjXaJf4gs5tDF6L
T4Nsrdb8uy3hlDeDxqi7WS6YaZz7kR+drxSPkoDmt1JxSxRr1rKMiv/Y+OLGKgjDqkLGXq9K5dkm
jXIjfY720UX7hljn1Eusme/JIllpFkrtw5Ulj0iutPT7aCH2KdXvV2gI7qAFeTa5eZ22pXkLUoSR
TqBhHNbeFjYBOjdxUnFFW7n2Qb4KJ9dffd+EJ98hH0HI0Qrn0PsdpSZGveH9PovrQ5bGFD2+QPnd
EhH2PlwroZcFx1b3bP239tpRkajq5Nvbybz97i2ubg4qK3seuJVRiz+qO4m0/DERqMsmC1tufpqh
x18TYZBv8+tEyK0+id7hXhSXQNqxtXY3LgH4xdxUxxIqjjlI8/l7JTXjxvbUD7vEGeN6JbDTq6ox
oVl5TiYeIz+5ZCze/nv5oxWk9sc5CB9GSxdRb+E1EJClctwPZQ8l+DfP2i3cLUsuG+M0D9dBm6il
3aAVWGKfxZSMtFSbVwBqE9N7AL9NdpOr3V3EI5lepRTvrQ8slnKGQNL2niaQOJZuZMpGA8Fno+h3
JbkChSK9q4Cbtd2u9yom+EPykP8uUygdY9iosqUzFetwFZk6kSZFb/1X1SHeURma02+4RhoCjtUW
RjkVh7ZaO/X39SvbRVHi9sTgiWnIsc6JYooMC92efsgPV7YMBg9TQBCnGPCeMP/55yEu49ZVJDJ0
Ws5xMDvDPvMXypr9O5XHW7GXLfNnyNB6PFFek5yF1toU04KJOLxuLs4dfua9lqrHuMWnymumxmx6
d1YhnU0x7R9n3+WtbfTBJkv25wndBPRwgsRp3D8Yp7GU9GbNAzZPnHOqV1yOQRN03BsBAYCnCT9f
zyvYlGWBMF0cfNgFTuQ6wVBv/Xo9S8GXTXyBCV++aN2yCff6bNfaaQKiI2of9Gbb1WDBG0ZFpiDH
yweZSxhsuoQ+e0AMdOf35wholh1fQaP9g1DV+SqHcQY90/UPbbXgpq0M1vmJukejFwh9KDGwzww0
ziP5mtncV73eszuRA8vHUfHxp+zwIp8G5iqL6kYYyux/JaPsYLFLk1vw2TfY0FoOnR8VvBnbf2Lz
sxiNXfEO0RRWBxFlZlmN8hTbnKNIu7MV3l/yvZqBG5BNHSM2bKijmGK7D4+eyjCBZ4VivgviFd5l
Xov3FXdks/lT6won097oh28/X45vT8u8D9sORTCuW1RHvhLIvuhnMneOw7+o3z9P/mKom0bJU1v1
fJ4/twHPrSFVy7GFS3RgVZXFpdMfFVk5HKWWrVzvvA0iJzg3EEqMHaMHCWORUfBVbur7S/H4385y
Rii2rDDDVlVwL3xKLxv7nqTizEinvUDoUcYaj6YeJ4aGn+znoMbHiAd/oO2jUkKxPxtUovFswutZ
UfVsNAJwoFtqM93IOehhek0J7scCEl2ZLA6b5SrW2DR2GRocoONv1HWjNdIUD0TumIYyleZ6mE6r
IroN03YvCl6+e3lCuwwIyhGz/wasJcsGipqqkO9Weg88dRNYUAwtPADXkL4PnamBxIypuDBMseeE
G/9Cx3M6NZVt/1uKxS48Kh3M4zptAp6Bl7yddY3owgUi3kEfTvHWLFWg5rnGGIwZsq6fbB93PYuv
svnK1YwktXiSahTe32DtCUpV6IK/qH9DuHwYN+ewiqu81tWR251sjLzOEt12e2o08c8tapXbleA2
gftNTf04nP4dA6frarpwYGxr6adlvsziOinHrQ1BFFAPn6ODl8N63cBb81q0RfSMEQq3YH4qS1Mx
C2kjAW1mA3sWP0atIi8bKHMFd3XiJInZ21nVhOfZicgrcTEMmKPGUjCKVtzz6uo0UfdtnmUwVguw
Cj9Ipo+523iDtwlwZtluyQGs75UgD6033gIyQU/RRqpjnKx01sT44B3OSDZ4oB/Lrw5C1bRcbT6u
olVOWbsHd9gjiq1FYk+AIQck4A7T6fydJJUaY7W8SXD/xMya9byuBLVmd87YLPRnFE6vimc/Tw7c
zRtGEl1HtD2iX1y6JQ46LVW6zGyLuR5e+JeY1kzg2leQsAzCmtdMw6yyab9Do6PS4XMOL9z/qnZo
KXvGW7cCwL9UHLwCK8GVsxaEZA+q572Z8CPDcZj1nnfEB2B9kKtN23NK1y9CwRnF6QwP2JEOp0X+
57rCEYLrGB0VtqiFh03+tCLd/p2mpo2zS13KlM7+hXXO23m6UFhKIaLaF6Q5rD+IsEKvl+QbSeT/
UXLn3TBqjK6KxfFGvJBYZIh/ThVMGgxftOCJr59TjppGdjGmVvlJw4iCfg9hPx7dHeFTn0D2m2Bx
zyqjVd7bc32Jj4jLsEyabLwk9gejTDekjT8caEnR/KooUcGXg+uUCFO+toP4XeqfLrDReVGbxDwa
Rl+7b9s2BPQQveup8NCTJeFnbxLPSOszD78tICV8g+FoPnQDKna3YjC+JlmwdlfLWPNHN9lP9H1x
ko4N7PNbbVr9fYDhSmEgik9utCPvQRBSUmI9swYM9WgDtC66axIjaKBIeM5+ZRoURGBBu8Rpyxqi
6kE4fmsLcQFmaNW8aEFu+PmR+5cJEkaGfiBaL7zjpMy/p3b48Lf69PK82snbJTTwaiPPtabns4D/
4LPy1A4YvShySbpfZcN5xgtzKMtHjknVshaTb3kZe/h15mjy3FRn9NuewMWyDUcfFVe4m7XHo0m9
ggLg+Xri0OazjLCMIVBmzFK0Ac6QyP7pAzmuusX5Qq8z/NGdYqx+FTb9sI3FVUE48TH6kHrEpzJ+
w67r4weH1lK06mN8NlCVRBA6j880c7YyieWrR/xzFbsvzq0fZBz1MycGnTj4RgRG0LOWcmLsrBE9
RB+Tam3n2UJ+D0N8kJPzPdktG7/en/0hxUMRu3Y4PU11HHBW/PmVPFM9TPo9pRCkk9wQe2WtCTOR
BALacOhRpjkRyJYYDml9kHoYOLJfSooMEmMCCZdTJjjOgak8Nw6jvjpkvveMy2eMjujyHEkP9OVu
rt2+zIialktb40gD1sYywQuafWzzPjMHDYrwkP6KoSo6cuNCIKSb8oS5SysZz9dEYrgjhCWIB/Va
pisclkSJb5rUa0swbLJSFOQpf/vxvw4aWZCYwAweN7CI1gdqhrNWKnF3AoHLk7OywiZ+PFx/yZ2i
I/Z0qtpeudhH3DqfhSBcFEyLNCzOiUb/VSF+Qhq77vo67m8r7fSw1TLqMT97wp2FLVk8NHDSyM/1
fNmXFNvFOmXHxd03WwPBdhrZRgt8CxQoTzN0OlROd86Iq1qwGC6QZysZ9GMamEEGoMJGsRF1tOln
YaaMkikFOa/qTpFiFlKL26N6kPJJhTHlYhENhBfZThSYW2s5hbZtMOjDsgdL5r5YzWk08g34peQX
YPDKsWWHLXj7z/iifCDq7EBQac3xe7htMwWRJL34gljTp0LWDEEEIUvJLSIWan2U0KhUJjE0Dc/e
LfZKKiJ/M2Q6/gstY2s7aDrlFaT1Sxmzlta+Do5+i+uXd80fRmlC7IhNAqbdZ97p4qo0anj8hzMg
VEYZY0IH/1wpxvvcF8dd0bDbzjBbmpaDJaGR8APmJRG5LF77crlCzpt4TyIvsgxaksRG/vKfV0L8
2+ZKQ4qwXt3Gc5cjRwZXJNG7GlrvXtiKVOnmvNBZhCpY7+uR9VAb1T3/ottbEZAqT45oV/hlybfX
cumCz7wfYvEsveQglkZpIztB0w/Iaiv/wTvWZUySBbEhQYkjg7EL9Oy1Bbzw5f3OK/5hIXO9BWHH
w6yQr2AzV8Y6ThUvghrN3zD0ocyy8QiNeX4KpPby2I5Lkz/iaWpNHvF6PuO+dJXckhDHc5ecUHUQ
cZ3KTV8TGBnw8oD84zogJQQkfY9J2SfxYWc5rux3Tu228ODjM+9ycGyJZB4hmCImGSNKjjNOoK8C
aOZ2xOFO0Gz9gGkV4SbWDgFOf9HeZxJCUdV1TK2Sa5wc/m/7mL1YlOFYaD5ukzvcYVvXgutqGu/I
wPpofoYt9hN5MqnzC+fUyNxfmSaVKkHiK8ve5ewHzPNV2Vx8jdk7yZKcAL887jcQ6HMIfcDf0+IR
pFmLx+LNKE4YPqJRW/SuWD65sZ1hTpQAinlW0cKVzMjJCToX3/4GicVNAmWgbTx0ofb28LK5OH1a
W58C28a/Fbpvm7lEzGWM8ejTlqGfISIaVlPO4M02qzxfkFKstqE6f0uUPvSgVcIr66r+hDNNYH7p
WWd1RrjI8yD4T9vBfWUCUt3r5McOEP5NlqPpaoCDezdO75Rvh3mY80wntjbTL6vuMYX1usyCDNfG
35UwuMBjytD1LW0YdmT2Il59MRXnjwjs8M58rv0C5JUvBiIbF5SUZb7db2ZpE+9bxuflrF2wQfxo
/eSc/twrU56tZo+eocEhDuJqqDBgKTMbfIHfxEsqpTjhO0iO8CdgJrI/hd9r6mip16PdkfJtppRF
v/uS8emO+BCur6ZO5Wgwpn2l+HZn1l/Xze6lsi2JpaHoNwmUO3GxuTei/BUNonjwoqsZqy92LUfr
XTDxDMPhMImgYUbvI6xoac37s71UNL4B3ysuD8qPxvjYKUZfLmxcIF+aCvMvwoyu2/w9KfYqQRqU
00EHyQZ3+SAT00LBwJE3n6q/NBUQ4vYBSGbFetPiomG4gNidzpUUYSKpGXxj2aVNKRXzbDPH9Q7I
MjSE773LQTg9XZpE0uFIDtLFfoQj/jXbNOC2RNqOrME/wkNaK4jkvV3TwcRL+WZwafjk9zyo6GJr
mBllVLsPJ9DelaGG0BWUMb65UAL6Eu5dFI7PD6AhGNggGqC+TWFrCRTyzs/Au6f0D3dr7JCIXKlZ
ZfUuZPCWi5GoLKflExB+5mWluTR3ThGqz6N0G1wyAawnPbThabcIpzQNa3ScOr/c4VfANsZjFVJo
pn6Gux694Wbsi3Uf5DyPp+eNEt9Zf9/jAma0yrPMY++tk99DY18gNFCP+OEJIA0zURwRrzglb3Zn
6sX78qMb+CCqk8SfExXWijxa8bzTQo6Uqox/fkfPDqY+uof7V4p56QzHDMek6Q+//sVBYclqVaFE
1sNY6yIjz2hBnmU9un60U7i3WrHYWdXLX/7WdmYcaDVtaDIJt8EQho+pjhSMjG2wKkF8/2joGwAJ
wOuO/5Qi/EhYHIzQQO+bASiCV59HQJC/Fp/lIZWsdi44HuAD+Xiz0NVU1PthG+2iSA9BkXwaNW/D
eyiycZllB/dZ1UVqIkn8hKMA98iJxHRRsF6DHsFDlV21M5qQMDMBKyAIKjSSPZOWPP37KgNpA2wY
NKjajbmIkE8ZMtuKIfnuKpd837SPHPaK7pc+iMhNPhoTb3qoUQ+Stvp0antmkEjrGXw8LKGPQHBJ
syvSxmBQ/PdIuzJ4W4EOtFUh14T9NCDO7chGC94foGxIKSfcS5IuydQGWvcrlTlzhA/LPku/5hZt
knhmpSpUv5yn57ZlP0VEtuqvO63zgW1Q4j9k1ZhWkWg/Iwl+wKarG76bA0Kdh8NikWLCZjeVk7TQ
CGFbiDXW8OaBUAyXg1DD9wFD7XxTKOumgxSy6YXDVXm1+WdFqDn+B1vG5AhOfGfzGDW+9YDEwuee
X12WsrWXpo7YzDIEux6NcPPeLG4MB90j9nhRHcwa18nmmHzK+G2mX1cRAJYilGNKB/6GYtTHxkpH
kOwKV5fFecfzVLIi9y66tmq3mbhdJH3GEurKXZCQN71ZHfCLaF1pcAl169moMapxHhEVOEnyEuik
neKJXcVuFTlvj2IG0i1mH/kbav0DdvZSaofvaOheQfgPZGhuJZ+1z5K42P2CGLqjJT+53ZhnUIYB
rY+TlsXNzBD1l0GL4HOzcIrqN1Y1vRNT42wS+S7vhDnMp9r6YDZfogGbO0fFU2RpHrVVmUiyg9Il
3t5/RH1VS1hUL/jWKnl7ymda3JaxK4dIu3H52PDYpp9Y5Vq6LAAaT/4zeQrXcOdsRvDky8BmtCTO
NQdgEW4GQpXYgwY3BxiYJ/stVN0euMk6GWnP8hxWhK9sIX+65n60VLXhFBS8q3/C6tW6PJrGdXSr
2s3vb/BetcOueg0+n/1EQbPvGoORGHFqHlmevYVQBoHmhXfrlFT5PpolvnVbEpIjVeVE1RfXG1Qq
olJ4bfNwXbUqRIirZpw4Gd2f/ik9T0FIp+Qv93ZPKed2bZx31ipdng6iZcQcBLXKqcKmFMO+C9P3
x9tZpNS9KC2XFT8xVnBathXa3d1cXutv24OIRSAfMeSPYJtgK81GrD+rC3cU/UExjchFchCmPNb4
bqLddJ57skHp98bjdldxx7HJQz0VfLIpZnnPPGS3oIq1fwxfFphr6gACuW4YfWPpeKTC5F6lV9ta
BOhmNdz/NW5FkcHzCOul5eXx9Bzx1hcxXPMx0KCl1VZP+VlV+FoY/pQZaYZNkdfa4tYBTu06KSZS
Pv2MKIHxyEm59pImSiN9ppIhyoZxw20iPBmvB666u6ZBxrvbkTbfAtgQOz6qTBemgQkxAX91npXz
UkIam9iHGho/uHRXJmj6fPq5POErz+kbbH4SO9Fqu/OCCmbQVJP6deB8rxVVPpAsn7Z4eULn64S/
s6v90c3UcBFVcXbs/WB3Sle6C22+Oobpscjo6as61TviBVkLMj9f+b1RuhNaS5hKiSWW+s2N51ij
mwdXSY5sASZXkGWoyghVn91arvvmPmzgW9Tf5zd/4d0YEFk+TRPTkXTnQ7dCui5OUEK/NSuYzpaN
3ZGrpetf9p9Yy6T+8RVj12ymve2hQH9VENnjff0Lgr3toKzLnkY4caY6IwF7K5ywaAztCyO2M32O
D2vqnmCjNSpOb45Z3vDQ8KS0ELKgdPOTyVnPVUTX5GcfZ8gSQaZXnt4DRMvFLWeUDh555Fb6H9Lu
aALHuVIdQMGhi2R7NEvilM9oFzZ9J8/bX6q40a0cKJVOP2QuzT0Rx2OlZufZyQt2w9bHEwOcFkLu
vJ10skKAQIUWh/KjmjV0Q4PIHR6eespDfWczAai+/foUoniEtHCfaCFetiA5LtTUbF+QSnF0uudC
M7kCf1AR2LxvTyoJoKZNFhkT9Imm2bilwdbkfmK3E043PF/nsJwcGp9cASM8nIVIeI0EIV38vDlc
1tHtxM9eZLGTSwBsmUxXu/ahuMkWgJDNvyd1YaHd0uzss+IP7YdEsGCNSOB66dg3nJhmScCGJM7l
8FcW4/USmOIn9nxeq8k1v8JSx2wz1OuDhAmj5TuabYpSGvNZmhfGEZD9DwEYOzaS5+UhES3jjzSG
eQAMUWJhPOkSs9YVbFMUPqykQcx6PiJI+Zm2Qcl1I/1ZQtVUlF699G3PN01rVu/GDIUPvI4Hr2Cl
G0XpATV39njfn5ryahS3e40ptxkz6KQbTl1NU3y2lCRadLJNYmfC80QcFlW19o6ojJGqRVJf5OGb
1oHCx/8yZv2f3+VKkJCCaM3cawhHL61/yJMvJFkX8R5+VBGqMgtLLZp4oJTlaR0E+6QkByUWVNwJ
8ykK/hDZnyfPIeQaLbMcpu/6a6atV34hWi85CEvZFU0ddgfSBde9mi+mHRGMIXMibwTxpZmomwH9
oLthjjmlVjzikhjHyLQJV6nQk7sGjnlmohtWGxzdjGBHZ6fED3dtCPIoUyVLZZ2VABSF6IQCvEi8
C6nc3Bmfuf6483NgllmsbmfCfveLvvo4Cmwic3cTnlMmYll5XONceARBdXLBUm3ZydNrI1nQkvth
604mwiPe0v2BXDV/32GNCV9V8wKwU+SJiUav+mGK5kEM0HcwCJ7ZN5l6XHUS432C4m++369YA7xM
cYPmN17UShy+OcItP+eMTP1mNOnnyWUGn5+hZWRfpjWsakrqCRAysBLrfWvqU9v+vjcP31GD3ZOb
j2m+QkkvSsT3p5sHfk2drGuM0LAzL5EiYzkWsBD/MODIWxlq+A/PnHvf8r3YgtAEYTNTEldUEgnY
NG+0mC5/i5oAas9mthpeQNtnPANR4Xb1roHtE4M8Zvm4NU4PH2RDX7+GGs2VVfZEtMlhRhEcgB4x
PojeseUXnrpyBMtqv1DhNAUfL/nzIwkOdFu90uxc/O4a3VnYVcoCwHXHCagmBHde4OSV9sMk4spX
022/gB7H6wtkEV3fq4jcl9T9WSwLSfNKmjOnXaB6fPZM0bXNaHMLuzymAa9UNUY4sU4XapWoQPBl
4n8XIdiWl6NSblJfAlKNobKxjKUGvVp7RINZoYopiEBv1dUrhWdjUJe5ZsC+zAISUu2ru7Qn6l1w
6aUnr+ztl+7i6jRTGwYifOYYDSgTsGaqM3FyOTjVtKMrx2zQHd4gyXvhFwlZl3NBGozH+zvsKlb3
APAWhtB/qFUeIUjSa3dPvAThDpNwSzEBXF/TXi24YqnNj0Du3KFScquzi5RohMHW+ezJVhe3ufNx
Qk3iybTW6UYXgwXUZH9D7HTW0IC2M3FjFb5nwpArpBiTGosTEc6lqVK3JhsCNInemIzACh6VssCS
GWTntYXnpP+BhGKQU5OtH996G8xPStnmAUU17q2C/mMLVj+7OgeRIw3kD8Tn+rQ5j1NeseT/H4vu
vR96RO7XS+RAiO4NDJl9CQbhALVNx6vjO0bueCgl+2Jbi0AMeytiobcMWNYgML+yiQJRFJ5t+M1b
Hhvazsb8XS3J/A8w0bzqah1X5LF1aneDYAFU+e+UErIr4yynL3jFH8b2c6rq68aRxebUctLA3Iu9
WdvQBPM4rgtbjkGB/bTewO4plF+NmsOa8n0cD+PHsyW3aTF6N12w8+bRK7iPbXGv39Pv0gPxBRg0
5VaiP+7hiWymzJ4z605frx9Jin4qfbngmFWvNKOtnxxO+1gOtqQ7qGSy8gK0YteneH0H190lQU1V
u16RaN8UZiRPr8TTZh6azNkUgohsmY5WuXBZ6NOkMv3GflxALexWgmBGFosBxrfjldNU2bpULKil
YcYBcCxOkOGgN+WNEuwAIzQgcfxKCv5ujBMP1F2TKKaNRAgYZdJngPN7eYt++19PJ1rSx5c71jqZ
E4XYx3s87AhYDMXoBEFoJ4rvu6fZh3lP1eLTdzPeal3/5TcU0B16fyKElcs+CYyTqWESx063XjJq
VJltnvGjVQ/VcCdIYCbsc74mVFCqyMUpWiO16YX0BQBkm01pjXqrLAryqKnc+MO8ztl+f7mmWXIe
pXBuGkBOehdHor/2SWkZ9ImJFVkCcBLYE5BZG57xXvRB2g2+Odov7j/hzCgi2wpvfTjxpLjq3mzn
P3VeSWfyQvnzc8G5JGu7aoiYfZ0c0pXcCG8FkimzBhNaygYCXE4GtymImjArtYfYxRg47Y9veYvk
qQdKKQoyG6A4RdSd/iHQKIbpHGbEp0q+VdCNS8eFgAY+gnQLOJMBrCGi5X5FtvfkDxjigGvWmL3b
iJnyPzmGND06hsJn6NZ+1tgz9rjtI5VOJD9en3WWDXXtD0woM9glnAbKv5Ro/ZkUA0d5mOfCd3JW
14qwxyFx8zqHeizfUx9uipgaKN7g/fOxfJKYzsAUHxisPGjEhwcK1CKDRBdXvA2K/0cEZHUUhSM8
BQ6EWTwMjM8ilSrLp+W5ra1ha5qwErfOut9/a0dKoog6IMW05rD/RPX8hD6rDlIwhasLBpOLt5oI
1/6ItiJpZXYUiqBLSlss9SV/bLChW1It4ms9EX6wI1FQcP3C3j/1G6jko+eALGrkpeTwwI5+iH8q
qKGKqJe9Fv4EjeEiK8IcBN9/mS6NBsbiJXSUaTOWe+WY/ucACyomx+BVwVoTpE1kUg3f/dlgCDaQ
+FUB9s6M6NpIQJ4nbXuQUkKh/+Aw1V17eueTxkxjxnvB/or5w6HvkWtHDd6KGOsC48rwxB/d1Oao
92Zbf5SHC6dqvv54EDSSqEkdqVHo5d7KPfFRFyXQsQn/fWq1RPufr9HiR1Q2G+Fgh420Fp8XC3yR
jX47xfXbuf2Mj7yieO4waayUXAsjmwjUk9/2/L1s+ZaLLREZCWbdU7S9rDoNJyRxSwJcs504iwEc
SQXhqXHPtLrangsWgxhz8F0ANhMOh5kb/tWCm2Hn8xKw4Z/jesEsGZtOUBIMihN/I5XbvmHY0A54
DZecrXNZ473H5XDXlw2NAufvtD/akJaIs5KpRBbbILBPYt55NidLMRg9Vods60p70Nq1RXMuk+EE
sjBw5D/LxuBZCBi3kIEZz/vObUnEyldD+1TPNu7r2AKxvpwXeETOmnaQhHlYzL38RBgJxQQOuRvN
Gv7YAR1V2/Yjp5kKu1YV/HqDSOL80KqnCbIcAHClG8CzTAMJAown6vKBEHk+2ozwJ9hh96dWEirP
Gj+HWF0RZklrXiql3U4w0sd9MgGDjP7Vm5llArwG35ASvfxj6WncUDwrJ+j7KtuTOJNvLAKUZxy5
boP/NZNwGysvFS0mECUL7Mnr2dBG21t15Rfhbyarj62YTlOm4EHNdC5HawF+Kd088wAneRz9aH7q
NSJhfHhg2SAjq2gOiEbZBq9M5s7jP8h1hYQwHIjnCzUFoGlwS0ZzCU75NgFDO+eDIxwc7nad1tuy
fLxuUev97jk9sanV3IO+ZbmwKeoFfDpfikML0SOE//N1Au+iJoENLi/cSS06reNKjiSxRNXhytL4
Qk3Cle1N8Wpbuat6J7C8D3hHgXwNqxQsj/ESnh8xGRupzsq7XA2o9p3bBLuhQ5aAuWI2HCASRQVZ
EfB9OiXWyHOPydpCFUYbMKyNJ8WCaiQsYWrWNkIoPriGXyahvCis2GjSAgozH7TGx4ydd5ldello
rTgd942kP0t4b/s59c4CXtvP46FnRfT8bfKcI0gPf1Z/Jhc+umgFMSv7JTSJodtZ94ODpiamQnKi
0KFukf5FrCR/gwQb7MPUbjpHJEevmxW5yD0HA9Fwf/e4boZdtzbjlHIolKIOJxemBE+AyXoVr0Ww
1krGnNqSQcGeJm2kixpNfr+sBhypuXkNXCu5WZC5/hzocesIJSZbdTEB6dSrwTHWNNq4r0O9lQ+q
LsqaoSF96ioWFEbDY4eetIVoGr9KFQCn2McTHDea4xBmD9djZ5EjAOcKMZ0zXfjphgQyIV5uiOVq
fIGNuxLaD7pBVPOJ+hI8D5k6/2MUtWGNMMlVUFnsmWKXPzf08hPhq8wW624rAFWNo8BoaS81rSfW
quY4QYaYyUHY96zOctOMZBV7I24/G8xdTCHOuZTepgnnxuKfP/1ZE4wo9s0AwIJBRI5xcTCoXVke
A2hoDybgJFfRg6DikH5KQDGRB4RAfkY7KUmWH73Q2Z8r8nxY5qPEPcBZT50ouH03Pqr7zjRFg1LQ
cChrF2cDsNDGt5Y6sDIaEHAFtJ0aLUnNLwlnfH2QwEatzNfHKMaQH+iOrUNjWDXPUlNh9ZSodY4Z
eWHm8WHECOZs/d6+Pxc6gNZF8UarJeR25a0yjF+8RdBNFoI9UmE1abdAfPcM6OiIv/Fw1AlF6fLJ
uWYeABcVnzfh9RZFZ17IkmDjjad3rPa6BGtlUrd1jLfF7g9BKkfz3HiM5EdQ1mHon1Y4dxazsQFC
Z1ZPsn7pzmSc1E58ucPgw7W/5a2uQ8JTZet8gLHZ9Qjk81eh4G2Pe++pzCg6mDzSCuUDYXdoeuDq
39OYbf+7g3s5kCPVk3toa7/y8vVSLCstn0zHfWGzAGq0pWhSYEWlJpTFkpzRdoicHRdq9TVENFFz
HHd2xFR/kIq1ZxXXawvN861dYrIgSzKZ3R/IJBvxv3Iay7cZRZTeSGXPWxpukgWDaUueKvaKL+KC
bAhflKoQCOHZ/Rhk98o8TWrg/vm8dFTvuEJA/FRmIYL+fdLIYtIgkelBwOIB9Db6aZEpR2NHgBul
S2j85aipnh7WjG5+cDCdl1YhXOjp0mkEqD7cEdru3eXoX1WPQbCIk037BEfxO3BjSL2R4NzS+663
6BimKjG3Y4qzgFM1eLye2ZK2iAuMOEFXuLecGgd5Zi1EzbMwfgoGWHtg6rRBQa5c07HmrRIwdBwT
9JrhsP+t8OvmWKXfmfQYxSWhHo/Z4+GZiaLrgvnsc5rKQ93OwMuZGVZpgxsKSf5tw4KC4g0b3evy
/BvwTb5N53wThScu2+uhNlAXEceNkwfpCNjOQXXeYD0/q8fiPmrwXYnw1yyphOj6LAq0A6Ay5n5f
QCSFa5xR8kyqIoJVjiQMlk8ClEQXUTTbniz1BE6Cqz6S0/Z18qZgg8q0KiKz7AY1Cd2mDJDHEcpd
xLDRaxXe7QaYvqsLSR0rz3QM8x1pLnu3JUIva3yq5WHrnP3pIjQygIX3hfrCBEfLmjfRO486dVzm
KX8LewI1O7z3lXZjCZtnRdWAgp/F+dPIV0lic7noqrNjavxiXplMK2BzBRqWMWwNSHe006kVQuf9
GbsipbXt6GYeoXvG7umcjTJmU0j0F/ZrHQxQ/8cgu+rp9Mp14o3ntxtUFyRq5BwCWH9Dt0/SZPHc
UhLJfHZU2nkbO547IPYLaoDRVq7E8joI1KQ0HedyfbLhNQnvIYwYK5yEGh4uORsrgE2lCfm0JKtc
EUv1Fh+royfr+/BSsc7gIY2lBugIdB9JB1dMSEk73Pa+uy1eIauj+OXHFXS5UNrGj86DaAYL/yWm
vgHvEqZegaZFgHUSWtsnbErSw/xnIN2o0NLWMI/OyXN0NsGw21V9wH6iVOdKUBdyCBXMxja+7+fY
Yg045g/OZzq2wzc47Pck5SDMJix4lvbojXjixh8/8f5MSvjgX/OKKESqL+i6vVkf04KuMqBWP4Uy
FYpYqBSv0ORX2nBPsUTVxMfM/hwJSrVgDtt/6c69i8D737jcYt5Hp8DkxTSinehZa7O4Zza9XzIn
UCRCKptfwYYa/ici7QTjYNCgqwMROraYI2ZdTk2Urjq60jkai3SGt+qa4M0s/C0YQ9baxMl6oFHz
tah/V5v/Den8KRU2qB/LMmQidMcobsTukoTK8nEfiw85GltRn1O9IyDbdOp5Ck3hLalbZZdgEqYU
SDyorn3efugUReFJfJ1NaVmPI7g3kMPfw6otkSWRypJACKZbqSuCiiplJ2450W9FfNHIA7/oHH02
rSjtUmN3pG+6jjFcyvYGIuVNZkOJ5bK8bIApWac0J6XnXxBc0LjYJ5ItFpUhIqjaNXtNNYMSB0PJ
YoU00U1rNocgaz4paGqYeXwL/6c8/CbEcIK1ssOH8mvDRCJsFpz3gunPsxsW0+j77EahdLV0hPAW
AV8OaAdFgcCokrAKSkSWQNmguu4ar2A0BMhBegSeIKz3iaj8OKOcL+xnfF7YDJ1Qlv1dUKrU6VnS
CI6fmZvceUakAsmIhh8G60jddWsQrRe5oQWjYjWjmLnn0YQrkTY7BUNmVdpBMyJ/0ot0k6CGpyf2
CciSoiC6nI196HOSlaB7wmDEnk0Inl06FvUOfOP14GMCGWk7K6Ge3SAUGZ29pLMezkXsARxDFPK3
YTkxpfkkqUkk0PUxAEjCUUNCKiWiFqYYNMzztMg2Xr1Mu9104nXmfQ7GEUeMV+tR1FgabXtozzHI
feEBGCuF1bTYtnYloK+EgNeq9Wpvfov0rJ2TfG4dlk62bYErZgm8pSSOqnv5kd+ekL/J/zGOc2D0
oUWafgtKd8GFD0fWDDs/Kinhm2U7JOO5ufZqXApyCtFb8bsTzlBJExYDxsX4pvujktb2loy83lfV
DNq71BC3KqeCgS+70l3AGbQh6r2Jzy6JePcpqdQ3EWe4gBI3ztD/1Z+aLCdDf7UbrEBY1EB6f9a/
muOitqpu6ldecFSZUE5WB8iV6I0jKQ/ZuOMePg1chhL6QSOLz0KvUHh+r4ax6dwhOZvg6ffaEgP1
Es4/nRw1+PPMFDZjE2MxoB3+FlBX9i73ntuic6ErHC/rmeRDiMGmprqo8wPdQhEUnxyMXSV5bB5v
K8HGQ11nrtVRgnNMqZ55yawQUm8Jp9pqcUfMkmjrIeeIOJmBiX29fTfPkaZLftZDynYSzrbJ3JRU
HO4YZyM5ys8DQghmtuFuwFcev1zsUK/n/kcFWT0JgNGWqfVPsrUjktbsTZBn6qBny3eZDtxGsspg
eopVlD4KKyOjxLx5Qtdc4WMYBCFoUCXHETUl+r7a28xQwMGxrFo+jbgqMG++Vz/hGKvoE0bwOzfw
+cUvNj0o5LTfytETqWGoC/lk6AjLVTO7FRc2NnfV7ODoqMcT6SBFQGo6yEFzMfqa4DJKWf7bBt/R
cyR9jLjtlyVtqfdOLpN/LQP5JYwgXU0Fm8x2Lwmt7xQYp/7ORHHBFPRJWKj2gLy7JdRp7r8F4Cm/
ss+RI/UhbSjIdVqG25ZH3B6rvjcBUJGot6FsXrPItarmDFRzTICHiIbbuBX0GGermovOFGdJ4Pd5
/op6+P/2lgy0Ff7THFBPqt+Zc0VfRTclJ8H7YfCpQ6jdgBjDeLBmwDRmUV9rYOChC7g0FSYqxt9W
uiZczzdyxC/WJaFcuVJv6Mi86afgmuV6oR32fA8mgiMlATFd+MRmh0sM0h/Yby5vzXyn1LPbPZJE
2i54blmYbygJyvbKK2WUuNQJ45BuAFYCjjKzB7JeVf71a3SaIbmaLe+kbpj7JtrIphSKPCQrvp+B
0z3THDKrrg3eqs3GroeRC0tWjqocz6pYCeb76zt4l4od74CUs32LACrENzDlA753SjbXgeUYFezJ
YAXrYv+jSfionXI1psIyOLCc1n3aUCjemVaz5RlN6R31daWXPYToKsfrRKA1K2uLgqT2G2Q2EbSC
Gtbbtuq1vK4VoEAxKH/CDiHsI0naxfO49OLpxRYBEBAQJ0waYkxSMEPWnnb17OUC6JSluoD0pgpJ
NY98FttT0/nqhTPW3JVZLHvIz40yXwOriR0q0En7NKU5Y3jsDcfKk/MuJXB1Tnk/GAs0yCJPCz+k
sGDYv9Py/y0ILlqejwMZT2XtwzFV2k3yJM+jGIS6GxyeRv/bAkWLYG6ZgbU5eJKh4vTqIXwzkRNC
sLXuuFdlPi4lD7vUUZLLkjUCeTJuEOxN9wCzEY4bsCah/DeRAnrqbh+gjxWXVByztSXLre7AWlQB
4B+XRvxeRusawiyOW/iGqtZ9FJiGhK4nsKyUnVTbuXmNaP8IryI70TgdZFPkJBE4z9H4GcR1j1CH
iYYYQeHauR8BNyANN146fcWHuPQL6IU94hnWPwVEzVEz0Roy3nZBfBggYnOHL1/ovrozaMRSPsoL
3/T805KNsQbgQy5qrNtkwMp0fRo0h6i5gX2BqwzgPuhW17swiaqJBaG0h3ySaKAPNWPYV66a03in
BDP/R/IZwrFRkOJhSrQDV4F83W5yd7Ot8VGjvctwsjfGgN1HbIzJx999WFeDAXvvNR26XJjO1IOQ
6nZ16pmn9nwPdviZg1WgwYYqX/b1AqX8diKkDt0yt0heXpiE/HlTu4GN7o+MTyygCndEOiS+BFIm
0TvV4L5Hnx87WjDst/rh/bKVML+cONMJ3QaK4ggocTpJC+HhAtAjzZoHWE4viUCAchKc3HgqbOOo
WX+qMi6wNQV8oANKjml2+7nY4BUBnZV/Ps0RIS6PSok8/PHaUDKOJSUCS48zWPSiNmfGe1AZ4n4s
ZMTzr8v9zOOVi5pwNvi1KGIhz8+DmPbllA2wICnImt0rNeGc30+aqgJytoPmNIf+wnLG7Xj35H7R
5aYSNZO4ss7EoNtsnReuvnljCdz+ch+x870koM7vACiWwMWjw2uMTq005jZIhqCVe22NYmjVmo9B
N2B25L6bay45O8kdKQVvfInAHww33q0uizi8whiWW2wkzo73xLMNgDBWSier9e/mIB5jfYbPP/Tk
8fklCoHYTi40k1Q/AzoJuo4f00AZESUWAL/y2MgD5/IKS38KdTJb8rF2DqQ4SvvETvulf2BKG99e
gWzPRB9nrL1YfhEr0vtKMU8AG3rWz7ZenSqNOTYAJv/inuS06Qe4X1lQ3npbt1veN17ni6vwrMDS
NtgY9mchBZi6SEOxS3rp7zqjzw3nA7ovnpSL2+62NgNOoFCHhq/8jPc90dZnbLIRTIRd9lU2/YEP
Ke2cUDikAoK4Nc+BFeohWpMlM5BikCWF1BOsxeTiCLsUSYW0wCbol/05WgTJFCOMni4Q0POUdhf+
FzgH7lilZ1SX91Gf1+2B40tYNwNKycLPwX77Ico+xFKysR0FgHCRA6/VOXf+zamq7JR1IQ/HSTFz
Gexo0GpqVgT0IQVzc3oA2XtOJCbY7IWfGnqVlJxs1GwiyE6LCLBKCGhMHsRHFTDBJBb0gGXBro9w
ymuT2Xf917hcN4Hs3JKnH2jnevATZNo9XhIeC3ICFFABmQasBgi9NLgxbR+iOUqxGC4bFIDniBy4
mDuv1SCQyhoolOQ5SIUi6tYRAP4xeTZBAXu7orG+jBXZpCvx9XOdA01qnXcpx4wCGV1n6R02fJRM
5FXQubEyFsLsNEw1mN+mXhB+gH32arEFmoN+JUvyTmsn30iEVUIhaB6I+jCUcPHEtztA2P62tDwL
8CqJpjYok946+AtcHUi6AiygRXPk85iGNWhqugniLFnwSYgIa0HpBkweecnma26gGL9O43o4Lemf
/BLteM4zp+2iNqBBGIgBOnpTgmDiAi/6sLXkkkw5C5R7hAQt0xGBT89xzZM60tDQ6C8YDeb/7DRS
gaMYy+GQU7G45ylApqHBuIpYqgEXe3Y31PSwnvDokG63jv7RkarnKeB19+QxA7TCh/VHRVFrpMin
PRFzkb7Px/MKca29yB7GoBS/5vjWeQQdUugEsB7GcTe8fTe5IrjUXBgeP4MrjWf7bWv23Um6GBwf
CuO08ohnjgj/WgtgT9hXqQpaOXqWcfpzwVJZcIpddQa4DPiDZmBoHxt2YOlqkyeeQ0ttXaAh3xM/
sBUQp7V3Kol7mqr60ngRENO5aDQLL+BlAz/1ebCobAnusk0vBxee/2GeWK3fN/JnoelwBXCLqMkg
k2UhrkjVHv5mdx7w0KDz2UPoGL46x57ga1NrD6wQFoPMDMxgoMact//Z89oZjkiMdVvz3SuvFoEl
bMOrJ9L5K8iLVgfck3VCvCoYGmADM//sRnB/sPdPu1cjACxKqhqyQMGUhtM5zbGWRu86oDfH485v
ZSzAlj3ftgOw5cMTSpTeNH5MgMOuPuyO4Ozgpfl304bRzPAYkVd6u9b9shcNUHuri5Ppz0oc2l0S
35y0nM1/N4acwFMd7Itzez1g504Wb2ygCAsENI5bDIUse+gySYpVtkIYz90aZArVjVRYchP6AE/H
5kghgY4Heotlea/O6xVrUFZ5u8t25VRq/aflsneja7CUN2nxkzlWGVzQbMYQstYXjY2yzHyWR5VI
erBjQ+GqkIaHhmEJ+OmelI8k0P0H9TI7Kmsga843Pms451IYMDczuHaH+zRgBcEQxyjjnxGaiMDh
XfYeem1GKM+Upu8RqllShSM9Aa8uglMOPGLb0uoz4ok6q7qm7nIaq/sbHkPpFp9Y8jQRdmeq2hFG
OKeLSOojJagMKG1Si8PhEDzo1r0j0Qwk3WAZl+IZuGnP92RSTfTHPGTP9F7n7DxhM92gDCcasojV
Yf1A6M/TcwaeIyWQuAU5GwTAAp+8JB/3B0AYieeZTOqYLsqRrp77MjiKazD88Yzk+gXNNjN4mTQJ
OEYXNbrJcRAQ1GlfddvOV2mWpx/5tNWVYm4frXVPZJeXmmXS4jSl/auP7dcjN/0iJS2TdB9fhP1T
tMjslvJTKJ+dXCXi2rrHCFGp3xL4o6vIfuIFU++YfBP9AjkhJnXVN5+yg5AxN0KARC+S5FJXxZob
EvLuL7rfSwR1wFBYevO+VWJ7ESiiBGb7EwPS8MUPgeG1lTmHnjuedlxMwamwdBteDDS9xdg7wISM
Ir0T3QtT6vzO0GmEYLu3s/ZSFMC9yui5hWGXqq0lGGUgARWw3sYD/RjOGwFE1GD2L0+XY76fGNYB
z9J4IJ30dGgt7ifdUYfGckxjuzTPCP75YI/Ok6F6ulc/MGqjN+m+pmDJ/Um3Qq+EA10/7Kj3txFD
HvfvWYLI5NljSbQAT4jCRAnOmmllhsFjU7w1bFhJ7NUo2+PXAwP/ccUtKqL6SJ3f1HQGBkiS39/l
p342v9qjWX+M5p1YRAr4I+xRpVZ1Ye1atEk+u6CY5BUoZtSu1VZJRmB2ywB+pa6L9bQo3ms3Iyej
CLqzttV8OGTxBdfRfniCWWYFbOhSe5QTQIpC5QHuLjPwCd7lECwnPSWfD4jeGORzw35nzjuhPNcz
55pbMA0CxdOTLb6ChEmwpijlCBYopwr3tv/M9j2XWyQ/fFkr6cPMkw0QoWkLLvsmHcpd9n6/Vq8T
1lcMCaPyPUHzLUbdH1jyY/D8yZ6lhRnYX9No9UHQ4hvQlCc9clk+EtU23tyl70jP08TCY63dudZ1
YK3NeCV43GnxwlMQ0yZNGTgM0/i1FVwUvo0NTxFXxfXPsyZxMJWfYcw14QkkM2MDnPbN5GuDoWCY
2Vqw7kzaTvMGl5LVwlPauMRIg8HHgzlO2PUqorI24vxERIZ6PgHWHfoaVFQWYTvGt9gixEp4OWHk
rqGlMxX4CMzlyWCueHT5xHTdij5wGFslHvR99v4KjMUWjJsIbMqvKLlp56H7iyyPHGKvyugzQOkc
xEBUrk9tt2WGmB6LdQBvJztuoG1el/y/iBQiHrkXNz6n0afhdEa1cVCEjRlC3BiOeQRW6bjFcPCH
+ZsL76baKgLm0WudFbUXijzqIK8/MqrSTwJ0x7ydA6WADsr2vfp3vnSR5IdTbTqherWrHXYtbLRZ
gZZ/p73fCKe80sG3LaYTQ4MF+N09msd4OwIeOPy45bK3Tqx0AjNEzUSg+yqaINvyMXnXAyYnIS9O
VwbnxZQhjBwMRvbOjm0xmfux4q4IgXgn1yyNT96g+GFxc6EeUi5XT6TNS5Rv8y8hHV0LWZoIr+pg
GQVi0YM68EgkBi6aMXrx+vT8vxGLVJqT+WAOtGzwNCfRD1jwnSC24kCijQCYyMiCypCAJDTri4bo
jWbhk8m1ZzPeeUx71qtCrkcA5w6XswTfQC1C9nrXWStVvj8Bg9nsgguGio9jifMYQoI+k9by3h91
kgKuN2JGbSXxX0R7CiiIntvVSUtF7RKOLUIbC8NXYC0t11mdfXR+iBI3lymoLuN8g27O8QDUwfjH
bRKmEEwkmPMO7nk4LrOmLKXUpGl5jVujgkmofqz/Y8OTWApJ0zFkLvqB7AvMyjLxtUmp3KvHjN1j
KVH8ccLCtVUf5mfKdZXFKKL9TrBc3RI5ffEHzliy1TbFaGChYgC8oEGFNGGicIc3HDrDcev8MO8j
pGYHuwshz3y3ZFBJEcOH0fndVP93vPRtHfX85ho+DgDIoXm1Rc8Di44321V63v0E3GFLAksHsP7c
cIxRqbTA1YC9ehADiDAzw4NV2Rv6OeAnBgpBi5Arnl5jLILPW8NUQhzvTxdu3/dOhV47yKPjJ8F8
bGZsDZQayyjmnG/oQCbVL4yxjDouatZ1HGZyCLIv3fK5hjKlBJJaw4YACVVbN66HNXI50el3elaB
PvqYCvuIHK4DbWKfn7+8QpYFB0PmdSJv7ms3yk5lILpuT9jAkETkkvpmCvGr22f0nCf5L8OwZmGU
9f7WrY2zrpAaNGIXpTIvyf47wQkr3A77IhjHdP/imosiMJC2oDKHRgaVRzLzwFGPDuxN+DFWxpAJ
csCyJU6qZ2YUPj2RTHgtl7nNLKgX/Ac0ODSkgriNfOc6H7nLN2Pn0O2X2sx6NUNp6CQ2Viw6Hpov
L5qOD9bFCeZhWQX5su582mrwG81BOk6XvEwBNiRXKHXT3MIAERJhJV8ZW8u1Pd8ltd5PbeZ/K3ag
cmHXRC9G76zw14RXaBYog28p78zFHtAha9Zz/1hcwGEbYb4EaLxhy3OBXbVHR1ZzGfuAyzdf3VbN
4tJnZq+AM2le7wAkiZtJlVoFIeKOPCd4JCsRvhPgjeRZkwbZNAP3DQDWtKeQ/uXQlTCC9z5kjHRd
dEO/g/gpMdj6GFfhbDjYKT4xMXbPc8lWI587gGH+5ej86C/og/tULI0QWkAuNE6trw0sQ6rre1dl
HcxWqw3YmcWOMtjH98J6HGEidFymoEua/Km27ML42Kg2PVJL1e1ThwLBBWDg1KTJamFC1rurAw69
zMBQiJYCr4F1xz5NaCJ+XPy8TK/hvqqopIqvoai+G3nLoG9ZFIxrpIDLnEIMe9o2AaYgNOUdamkZ
0z0p+awxx3kSX6eLkW2DJbZdxtcVpWA0CoXKL4XLYN8VZfJHKmpgRfzP8/EH4PsGrG99UsCoPAp2
GWHI94uWlBOHDKJhOVwVv+X0H+TzdhYsJ80f6XkxkSry+gsNDlZ8pomyTORbODd4xtDLL08mjTX8
/iw2FXemio9ue7yo+CuwpBru8dBw6SZxNgFre9tPwIpvNinNkD2oQ/KcLwJPVxQkwdcY1IMBcUOq
VUdpV5Wc39ln85jdtwRV63dMDn+iXzROPnnPHRxQqtOjNSw9a1PKij0evs3PtFZygXn0o6t0M8Yk
hkzaI0LJlVCRElE9IrftW1iDcs+WOgTqFIzOv0FwfxKoMiSijBBbOa4qUIthFvGyCnMiNZMM8ftQ
0vfhg/lkvEL0NZ/At4qaKkcfU+1MpemtFFbtA6IKRYrAUEPsAO3Ser/rtFjhex6FP8zoR7K0iegy
MdXr3URkRgjo8kZLgdVYOBmVLwR40KGr4pdFv/tDuEvcDb1+bqgCEO584h0dUOmt9zxZVwiXoSIx
atUxdFlh6ITWc8+yXAMHmHVMHT/7kqnRfhjkOLw4ut/8/XsL9K2cPXR6ga9P15QKqtDJbNK5uoE+
RG9CCggMXdOfReflkUWeq37UeJwA8Iq/ht+9+7SIbCeNY5DWZ0E75gF8EtnxgEg+EtPf0tBMNLzK
4LyLCR6wc5vDn7spyajKYbxgUAZCBZRFF+Zk6uXU3VGZ+fdPQ/QtOsB3KvsjYzY58CP0vV/uD+K+
rMZTZWqVbRJSF4/KWtvGzJqIC7twPNLMsgD61wdAHtf3H451k6dg+LinwdEszYqXzuj5I+vNVa41
hdH5J3wRVpHj+/fCr3LCrwC5eWNNa1y1G18Gfy1EneNtj7P+LcTwa4uAip2q+05eGYIvr375tb21
ysW4uIphz/XOx1tgnj6Xe2uhX8IOXIs4/JInCaLRtgHAoiceNMRv2KcrCG+LkfGz0n0E8N/LpnEu
DnbNgHYSelSfudDHMKDJX96ZacjQqdVrWJyEQguAh33izj8MmLA6o/Is1Kj3cvs2sAtKemsL1OWM
xlf+vOj6j1/DjQH0+X4vWreyPG3SF01H+cApe7daZhvo3BELATDVM9vlBzQ/TyXZZAm1+TTyOS7N
XILGBMB34do6Kq/kFBmrJW1hv1iIuVHIDrtTxDGwDnjry9vFiB4n8lIeBSO2GcXMu0Oz0IhcEfPJ
UxWLHt5o2VVbhZ/Bei38q+BEe5tf4+jsRd1L/jz009ehW0vnciDJWm3J0L1cGIi4MxTqWBAjSFoU
eRVmFAaKKB9XGVLW6LXq2p0Y0miFPe42G+auX0Z1+6+pNiD2amktLz+zvzjw1enyRxgllnP6YGJJ
yMxRH5OL39oKWtSlHDzIRy+THiQG4iW1PYnb9ewrQnnCD+c+GqWBcSxvbEk3ibqWqBaIC3xqNl+Y
RRsXALw64np3bNiJRjEHAe7QY+PVkCsxhkeRKG+oEF5X3oplt0BsP3qxG1DiWo5IIUonSRAihs26
od/aRGRfCsCJSL7q6v0JFBJOGtyE78i2uvhU4RyvENV4N4lko+3JJf6JCxXt1lMpDVrCjN6trqSJ
95ZpOPrKaNRZJwO76HpOgGw/8tf/ZCPHDEqu+IY8rEDV8643sOjjnPlUlRHPfoTaZloBw1phjSHJ
pGMKytAtsSlIW+S8y8amiiolHuBoj3hTU0gxSTeYRj4TBv/p+vMKJKVS7fO7xDJKQ3rW5qYzIWhn
x/DQYdOaHpbJXrSD6zkv9lHC8cpbymRTuX5ATjAKJxKEs/1cKf5I5YzGGcZvQOu87oX+aGQNRre0
H4isjeKdm6umB8+dN16GLTODb/qj4s85bo2hJLJJmHfHW0KKZgRfqscVnWaX4UU9+V3kcZoy6Lj7
srGkCvmpGITT7OWA2pqdwfzmDVRNv+MmTfXaZ4uKNP55BAwiDRqQ/4P5c5xJ++epPYaqZFT32n38
a6jE2HvSjpX03N8v+v2CbllNc5S9gTWFJzQQFpXOjLzOo7qD9dsZqkMPROL7h94j8jjzcFJ+11vC
fFVM/GTzm0PpWji743UkkrsO6gf7C98cYmnH6Jbk/c5Q88Yir1K4aTLyG6Jy8To0cnw+8jMpBuBe
DwgYiOyApTpXifvfXjTwMsR7BpkzRvwCigmRmv9Cop/ckXaTMrpf6wlpiRcX7aiISt6NGiUhk37M
wjdtUjkDhRSFnV6MgP/mvohB2gOCXgMEz6MhGAliOJiEKV/Sfc2yESEvMM6IkPqukqTFI6RlHS9M
wL4Ybg/ayafIUcVW6uyyGzm1MwZQrG72A80/hLGuZyv3neeq1vjSTCj4VueOCcCcDuEDKBEJ5XfB
0BEQJpKZ9A1woBl3mZEr9141nblr+Q2VzCvVDdB/L39rAkmA5NpRlsKxBqHJp7G+LjfBOxpiAmgc
VxZwKgMbF9B3pPGTAik1sAgpRjXFWIXR3fV/XnSYLgirsv1WQ38SFoEE5ZK5jn8ugJKE31tW74DY
wngujoiQmpFPYjtNDwo3o254SXg1cA1BqkvyttCBBItJFp+FH1zeFLYiAZd06adJTfQ6ZVSDr4no
5fkFz/V2J87RFgN5Z4Gpqcs2Nj8GObuM4k7cDW2I8SyDvJ0Ka2hlDUWfCHr9e3YvyQAt0BVR68pT
TtVqqVEQdLAlkN43z7yNZmi+7k76qlOQl/IaVetxRZm5Xjku71G0vEm9nkM/AFd+sTLnxBKc+Qyb
uzk5PUy6WDCDlPD22q4FWGzZMHMBKaF73G5UMqzwg0BU2lZE5A/zDt+xhmuC2kUyGsoQa1zputzJ
8YdG//iVWkAunb6JbXDpns7B2T12M6pIy4GuDz8gp6A9NgfLGPvWQIlPQ85c+5ChXx7RQuZHVkZe
MTv7lfQ4e5k7giQ03rPH/7VAygY4z5trYKSvx5y67Jy58/iyx1lMuwjfltAdSgznI46vbFVYVp5d
t/lHvbYdcsjcgI2UbPSAo8rIFQEIaBcVvtrwQ9Khl0Bf6A7QPjw93y9SuKmHl0c34s/EVsCOm8+I
ArBiDs5esnmhUfO1QnZLyRwD4sBT+5QWCHHkJbr9Ub52tIya3yS+I95bFeN3VixrtWGpH88msOYq
xovvBg2WX00BtoMwUEFkfdEmEnTAlsR7y6XL1zZSviB6fCcT9mcjdoEItG5PE6je/Jx1HncmUMzM
rPDfSfhSMMPIhK5faa0O6bmGaEaFKvfS/wlT8ew/LiNqnbYQj37hu5pyFXsTYYxgEIAqApFhdJk/
B/R/XxXU7pMrJGvVbn9jYmNBumWAbgxe1DN/FM2hYi5zlga1PQGVYZQM0OH5Bsxu4EeNEWLzdIeC
qHZocfPdKKHOR4fSR+GGgXcXXpdEBBiB4qSM/wTMUe44AtemzCQEkPpKGhw3fmFe/ZPRWrss5bHQ
WEw+PSfMw9uDl77kM8qaNOveYgF/PQMf1b9+ZEzXCTAKUWvHLgCaMwcQ+WQFzZ7vckMZD/oOQJPj
R51J+xE/EBrLH9AUUWY4QUkHh12ieSpZVk/LWQ7y5y3i96jGrMsQ6Ni+s6BXC5KBD1qaRI0qnmyt
TuMBDBrG4bM/OD+TC9lpNRkAwON7jGKjTYkzkfZh/2QDF60wkicmlYahv6LXnLg/R11ShE8vCxKA
Xnx3SMN+l9aew1ydcjU+Jth1wrVw0O50Uks3EFCKxKA5v1tPl+yVw3e4eXdCiJ3UDtDZKc73rZtY
BhirrNhYyvnkKTtNFKAOU0qlg9aaSqjgJ1nI9jMqHHt0DqO4E2P3fUKpnMN9+lsWwHHiesIc6MhS
snCiGMB/bcp5lLvBSIiT7W1I0Y5lUNHZYr5PkAjD6BK4jPAQ1g0GMeodCbiOEsLL8r65jjPuT0Uc
b8hXBmh45O8hQ+euExZoj21IK6LdNDD0Qi59izF2m+2O9PFJn1BxCnumKcdFqFNSQB/J/CEZ6YX1
UbtDEqzCUcH4RbIQGS+NBKi2XdfJ6BNviXcuVEWrbob/sXsG63T6B0Sh6yG+/7BG1wzsbk1/yZM3
B9E52f3FS+HHZ8RiVWwdSwuszEMjeOenJYFG3ncnYWOe71/D22eRxxWDdU5eccpMR+8LGJ5q5IXN
2KJ9kmaHYOTA1ncw2/Mp8QJZC0X7barJTSSErRYBHR5F++Vs4AhX3ClnON/uAE3yM1RxXIXQGVJv
xxrlWaZM5inxI9sSc8icbCVV8lwxbBcG/nZFUgubexabOw2HIF5P/2QNCbKhnePSbiCptIPw4fOV
9ekqKwnWPIlrJwyNQUkoIQshmDPc8Og8FL/U4aR74WdK6+ZjF2i6TlD/2xVYr1XI2hxoczEQE3k3
aJOv3LRJ/KYm+MlPD8UR9m6V4nrY81bhgV3easBU/IDHbFSfKnYI9DMUUe3F4sAVt87Lm0j2x2XM
xdPWbzcW2OnHT6dIUV0aATDu4Ygj5HNtlRjsKcyZEO0g/0TzMNzNiV7l8+hdXBnrbSbhFQ4zvclP
+/ldajA4nUw1pT+fB3uzuQTcb8L8lvnl9bpIPqkeLzetOgD0y59iGUrxYm5/lhrqODjuje/6x0Ce
Ahxmqaj2zu27pWJ5UfrGhwgE9miYL0uLpmmt1Q02/wU0vuLzwb9p05tXqmXwEM6If9sgLyOCDFNS
GCEgvEtlHiRsrubkVy0shSOk+Csu3+C2oQ8W6x7b0NDKRrcx157APB5uarVpRRPxfqvz8Cwb84Rk
uTnPMXVoDzhmLShe5uhsxWYty8vgqXZLNl5q/nt4Nn0X5MpBbtKizBtcI7o+npWMAeP2c8M6Ovi9
vAuSXssvLMlIPCFxBA207YFLyBZQiUXP8iW8BeeCmH51+wv4ALEXcilkjo2upRnnR8PDOkbIn17G
sboVl54GkYNU7RKa+PcBcjkKWuU0CC3YvRhgLvjn1ZphuamwkZZMLA2ue0DXPfzJJ0RFQf+c/y/2
fsLmsRP+1J2ewP4otiAGlpXq7tFmroNmJ91EsYmCsUh9LppQQV9/Xhg5O8qLXNYNlzhdQlf19dXA
aR51xs+ZrPmW/o4Kh1p+a5HA9fYeFyJLt+qOZ1FeK2fgUwT7ABTmU8OD9WkECG4oiw9/XtIA5R/e
6TUIebwvyZDcMoW4Pb6a/MClLG+p9tUS/BoG044EgfkJEb5+3+CH5FpCL4bYRUqNUX53HL6xcPc5
5B9KBFLQDhDx91eV1eEX8bpSPAfv1GAKyrGnl10IDPVNIFZ9nERDPteGYVvJg9mrEphGgsoh7rGO
sU10lJ524wFewQHrtt3NqaD2vrvgFs9qiikR3At+18ghVKz/hvUHEwdGCrjIb6euYkkQZgsCtNNq
mVqcv9PfxRbkrxgO7Fow7P72P1VgIQsLp3Z+FzwqNhc6+F3yAEdLO6hvtY8oQGxS+59u/t/nVfiA
MTr+HwHyRrGwb3rgLz7+pkzDB0aJCIT2y9+zw3HchzcCVwJuldSQYwRdtXoKNVGPpWL6AoU5LOlH
Ee+xKdkbH75VEalmDyq5dP7kSQOIVVNoQ3R/8/Do18cqXtkCxajbEW2YSxAS5tkb+18iWbIE4V9N
Ap/8ZHwOyAaBGoFZ7pucECVbS/t5FKlJFsVLASYHaki6x/OhMqxQYz8v0jpq3EO4CYDdqr6Fu4ee
rbDz8z7Gn4JwdQnSndWU0oAMbGCzAbbX8CA8kDgKluFYN+8XR/rsJpzluI6+amEL2PrwLZb9Rwsj
kCFqPckNuY3SGBItBRgVR4fJ9haFOqX6smTm5DMrBOUsiC3QlWxYXTCoP9CEgq6b2nyobvVDEtZh
K6QzBTxhBI4Uh3qiUKykTPjc3wiB4CVUJukuMB9pFI7zovog+hQB6RWMs+GMKqqCTnitdG5iOdic
tgT+Ltk7zAg8bNjJulM2t2ONJmqyFOeI65EBcEfq/PGFR92mkzg7sBWVBnu+gPbwVy1wuYKsLwIN
HBx6T+ONvTzDu1k+UteizmN22uydqWZYXaq7qydsO1t/ckHwhy35XEZR8UfEFyxZfPgMRlkltWO6
nMoiSg4GQAbp1VZOsZeWnH3U5nYxo3UgOtUwelOXlVijuAZms/EF/5068rMpiZWl8bmfKnjmFAjy
do28il2PzJK0rgF+v1qllVmGXmnvGuDruIH2FxAfQ6apoG1fRqa3tgxA4TilfDZ2GJas6TfA8mBt
JMx08HNeDuKkYo7EAR0pdBCsn/Fkv6Q+/Qh6QQ+lQ5xHgSDXdeuVDYo8fX/5qDoWRZKu3+SnF8u0
nalg4NIUAViqQTJTXoNo4nl7nGX8uaNcU6RAZEqvsq4STZwoZfqBMlLsAaHtLHCrJ36Mm56+bvho
QJyNOo0LlRet7yY6Sq/l9RMWkhSWOhfbY0Nv3CjpI/Eicoda/psUSK+tenTOYeMeeGfREwQyf16h
y/rPs0P0rIbpzkhqE2Z/BWnAN7VjoceNDmhbnPSZ8Aw0qAUEYFvjr/aX68w22hxCbUYjQOVbg/bY
4trwcCo5ggZd8gW8IpGsq1S2kQhnLCQ7aPVKhNl0h+5xwCobQMWEMpPqpzm2v7c44GzmkhYAyVA6
W+5OPAQNoXKFVsSHcmtuTf3C/2a+eaYgQ0WZyqRbgc1tYzoLOw/Ihyun6JlOo36WSeqcmhYbH1hC
W43C60231z4FWTqAVAB/E7v9O1eWMw4UdLEEV2IdeUh71MjQ+jyCtogBKndf6PYZQ3hjeL0Zmg7n
tMqjsAivzltXbrQmsfnCc2fJhWE++97aK1cRhnKY5fYZXxfReRF/yRQfnInlRURG8yLq8Qd0haOT
/xw1ev1pY/iAYfVQIc1IzgTcE5pFXhRjGeL9vgPEhtxGpylY/RrZQuVVEuWZcZr0ChiLs649oJRf
xY1AyBwrArioyFHnMVhLJfYCgBN1TfIx6yKW8PMF30K4bRaItHgu9CZxIrkSSfWIdSgxLVAGMdrQ
gsCgFHyottJ5VBH2J3BkPerM0d9ZbR+fOvaCyWu8unUwmJJ41Tt0TKxed+9+Try8EkZKpdj7L6Mh
hHruAb0AYVxl4rh8LO1DB9QNmpqNZ3YRZCKVZJYVVVludkVEK+PeZfp8xSjBXYEZEwLy9pZNRNHl
xuh/XVv2Uvr+ow5DzVvvMigSUkUwZFEmzXJ1xxRh7VWxS9GlTRz5LQfDCqxv83DQb+1HwGbfWgQT
I6nEFn4k3CkYT/8wFFkOoYJfH+99bVMh2Q6z0plCQaHpaNSepS3CwGpzeAtlMllu8IXa+Oo3gA9N
UUOm08DCX7EjOWl88qKsgM6Zy6adEfqadkPlsK/8eNzL15PdJLjtIJruPneDqKk5AY7L1zvdyNcq
iItoqWOcwUmRlaS8NUvUPQvkcDMP17IZQ2ublgmtxvODNZmgNc33uUVj5iHtWjc27TemTq96OWt0
qZxq6DZJQ+8sbhRb8p3XU5Qo0A6GW2F3OxEwak3otZ1Tkuni/P0guPQFBSYEH425RYTKblI65/fJ
ojXNR7otj4HUGzRH/BpMfManR+gUWmTZriNDKyCT9w8SH8BRrSchcJBG/jG4SEBeKaMBxVtHfbSk
TgbaMeN39tySpFbhOBjD+59Jv8IBlYdyDZx64YwmNEp0uoesS9sb0BeK66+8iAbKbb1IgGJPTdTE
5tRY2kvDRn38NudUT4XxczB1BryHUd9l24208G7X480xn7R2tZhZbBcJcCwVrYLCSpVuz/AQkey6
MYtDprxeW4CtRia0oYsXSA0aCP0G/nA7IFcerFBuS3YKgORj44CgS+X8eFnOr+WX8DMrD4eg8iqQ
7YJcXPk958xFGv5BeURPfr5q/yf7fTWK+xbRYb99kpCxtR5/7CUJDeDOSV5rP9awbrbW4iZPEo++
VX0eb2s7dDQdjpAJ1ABhq03P33g4YjlbjQ3rzQYbyxeaR8jAk44Y/Q+F/viWr4AYTHwbdo909Q9y
IOUWNky1KJX1QZ9njfSFm11Vjdl/8+tCYHQEx4WTUu+BzwadDRX3hWlD4g7FE0GDvCCAMtIyhARd
QQztM1NwSZaNJngBVtNeN1CqXG/5jdbG3al1vioqN0/XhWIyaGUrLcr/LliDHRIkMnUM4sQMRijX
H8n/vcdXTcMzX1xb3H+bLEy/0ph9kbvLKNKhG3cYo5H7+2zgQ8vz7Uqz30gxjJZ52/c80zcEXthM
GmpuJsI+KbUMvjZqUkKVURhKcm1uvtG0TuSJ0YTKUySo1XJ8JlJF2CmAnyjkFNEgOFJHAj1KOcnM
pn6m8PbZnIigH7x2fHVOb+IGCzj3rafLu3e5YIbZlUWE22QgftVZAHBf89KgsaAAzQO/7nspZvPB
61AIrPEY7SlHsyd5w3ZzUMUV6z+RPMtKlJd3toLfdTDsiT8VYReTULt7QcuMUAu3VfxCdipltH7p
5Q//OnzNZc/QYP0w8vnvPXmhKEiFbsHONQtTbjax+WF+dMzhqhIvkX7DdcihtlD/baMjWlM/2I69
P6DqDV/KPpNq1SUKhnxAsevIoTNVarnmQg++idmVUzIfZu65rQIZHeLwyO7g2ul/iLgmNBecpCoQ
IrWlxS3ffyZyLR4da+ex04CnjnA+sM8Ru0IX1C+DFYNuJR7E3bA4TxuNQ19x/myz3YZiscTjJzcV
l1XZftBZtG+eJ/wqtYknd/B8mhbFhIxwOOT8I71C0zzJ1FMTLY4XuWubMS8WA5DZHMwQWIksItvf
pHEirR0GuAqbZ8bVgZeaZYhH2dy5z+y/JN8IZxJri5hh7DwkL4IYHx/zyp9+uAe5Xre2siiuFPE3
qTpyRruPnulG3X7elh+gSJ0j9tUEKR93kxQp7+yyu7Ksm49+n7Anjipd4v78AZiQrbF2PQeC3wQr
i8+nl5VRMJ67PI1thvgF6c5OXJz/d6a56bJ1X1Le7/dZ8NFfeFMPAWw9RyB72wX3Y9bCEFF0PVGm
C/x6HCemRJa6Tdw38S1IOMvaRQ+WG0BKfjvdXMeRh6FQdvZneFLkvHUA/jmqO4VzIRctGM4YK/46
95Gr9Ucq0yeTaaREmpE6wQtwTuhnqTtQM026Y8UMpCaLZGYMLbgSBrBrwKBCa6bNt9sJOb0y3P1D
9EtZkp8GNttpwzhZSN1BOYrVzsVOLhAJM6qGWfWf/66UeVZL1qkrAT5e1BrgL/IFOimhr94awIS0
KIQ7kr7SPCqfKvJWBRAWT/Rhcg80QPgPMPC9lI29bTt4jcC+ckK8bnMzoO+wDDtVDGvnoNmFqbtV
/+2mUmsI3YikFoXIxVpzptKHFBUk4DYYGmACUoY7TMUi5j0W7cw/K7+KHooqQZ8t5ojpn7PVxkZX
a7n69QVF/YYhyUpQSwmLRqlUXs9n5EscqbMUr/Z80SyhEnnYaPFMkvNNbDN9U1Nydj4tMbp32sXG
qqKxhsvH2PXNRdf/d4+YOuYX7nxYz07W0NavLJPsgDFVwzk8RWg1xXW5JuGUo/PxzUco58Y45eHR
Z2z4uZJLKC9oSMZkgbOD0xdH5qfcJAbts14tnlcRuADrYNvHMmI7ltNaOnJkO5+CHM9OJLgXyqK/
/pTcCzpRhgsYXuJIlaRSySPwFGg/mBwwysEuvLfh4hHzU3+maEBC5mf3EuB2dtm8Q3Sql05ipeWl
aCJP+h1Q/1CBASSX2ueATqBjH5u7uObegZsemKcQkH7jsHgSdzuuCwjI0fWBnAXlWRgCJwQCMSE5
mRU9JoPWaLQsCE+JrC+ngV3I07D9IOqTC09lqS9HP6LPf6GLiFzDZLhNA4692Mp3FNOuto0u8Is3
GAjfjoqeCzGEHxwfM65c/cKc64ycU23KapBuypV8pTxgnWkvF2pX4zZw9IaIk8xiRHfBR840euLV
qLNZ3Ut2AHlS33Fk1j8YyXs+eX/0X4mK489jlmdjTyHVS+tRMzuXCdiIJp45lTEYDgYLMkO5/7f8
AlO03RRdzBgGuWgt8JB8RsoZq7vSxfdmaGpCF6SfMs965AkFfuVi6IY8GNUVzPkWf6j5qaqxn3AC
pbm4cchiVOiENFfup6w1nRSPqm91chTVZME6wLKsagg6LpORWMfVU0DBOoG5y2bPfB4ZDgP9u9C5
68gB09DJ/eNgU6BLSGrSGc5abcZq93KqhayeasLv9EWZ/QULNDvHrxPuLdE3Ki4AXnkK6/oVZfqt
Z7Y+PD8Pwxlb6yPjKa7R5Z7FUlKWjZl9U/58FCYFBtNOJ/7WQG6zIRMXyVFjpECwZ7TrHvaO5zJF
sf4n8Hdd91CxGhniixv7lAxgTj5rXPJ9NxYSHnl8EJkg+SUYPSNQVgkzpCwfw2wGzaHZy/OYIc3N
YPGruPF8AlrLcDY0wMD1izSGUEnoOQqGOxQLYe7W1osP/TPOVnPR1t0G/CSS7z5lQxXQSQ5eP4o6
ZsdPsTL15jlEyzrOM5He4Pa7SnVxO4hOX+7SKe/eaBy3j0pLCXIaKrg73AKi9pufSe6rq9lEm3sT
4Omu/t1AChm6MxBib2prJq2UBSfQdJ17s0Dvz9uV94QGtznwj/Hf+A6WqdDh4Nm1n8Jucm7h4Pmm
CIY89+5YDR4aVuXL+F5mJLMNytU60y7Dm9s1rLQpLPlDP5yUsntAP0saJ00CoFXKlxS4jkPlSN9L
hmLcIAZsSPXdPdgIA+v3kKm8h15Jhhu8N0xDJIzDxWqzl2RoPbVnyLTjREYM6ffogFDcTBBjLW7O
pp/Gwecgp/yK2nna+5oTIAV84RLn0jbDK1e3SAj83ciUNTKp00YLmGzGn28Z60CwzJbpXNbtLHsc
9YDl0pomkUUgs6VBB7sGv90D2QJMI0ZE67R7u5B74j+1qhXd5/i9uLsUuy5z5/tHOQOknb6FrsA2
MYRg5A+eXCvUV9eL4SO/fEK/CIqYUYPMEUpTyiI142OoTZviWImVMAQIYyq+Ony598dJ1PiPnsY/
AH/h0A29yqvMUrxFeT+Gwz74GrSa0c4m4/FW9+qMaTDIB5XsTrlZoiInKRvLu+qC3KDQHhE6nwGM
Wsm/WgTkkdYCY8vXjGipV0E1nZ/3XsgmD138IMK+J/wExbEp0Md+5TpwkqogQq8B+bwh7FyGetqx
l+VRbi/pERLtuaoGLgbfGG2Ot7RkWOxkBh6MBmRpg5bult7kOFsT3SJYZbh73TV6Iv2u0MtDHxUt
Ag1Fea9neFVoMZptWJYarr/52J5eC9SlRqoxElddTQpNUKLM33bP2onIMgmi8QpgcBm9u4CWmabm
mwezRjZkfxCkLYkCtZtvVcCxNQHIIk3WRSL2s0eiFEmVCZmLfzcz31MUWRhkTMx0Vl1LO4Z7eZ/a
QG0BkhKDC9KeFbn8f8Kf0S2d46SowjUA4+rkgvH4F51E6FxeNv8+JujGy5eUvvIIOctG+kduYkbB
r7FHmWheRxZ2XFINqIlHCMOtRYSh1511b+25LtzhcRWcOg8AnL2n1KGBV1n4NcAsC7yYtSGWQ24N
dEmy+BR3Lw4ENg/92Na4VTtCjjSNYrMqxz7m0fx8SV29Ey373GdniEAqQs9jLeIPJxPKRo08HrrL
GBJ0vH3Yts8m53csyVxhsV3Nsz7TINCcKVuDtQf913vNFfkwPqWvDOeUQEPRSbtNnrMa67rfMc1c
62VGsp5kBmAy1Nhdc60kmkblCNKoJrPuZzvJGtyP+7DQAHBp9PFSYCZs0CwP7b0nDJYRk2Gc0ImT
JUzg673kuF+uvMHyDQRNTCjmIVgQ4m2evwGh7pLs4ED5lLVeSVg8EK3KfZ3lUJzto+a8o4yVBY8N
0SYPPIWZ48yWjceDCcLIpqRukzoqVRq8szHHQi8hDjUNR5VNps0MGjt5aPzThd+vnuY7ZpsxbO+o
/3uXaX/FDvwL+CWOO+yTLLHKku+hvKI643ior0Q8AbUZ2wiiPv2zk1pO4uXlaIuLH4rjStUENroT
6uzcy93v87PW9tVVLj64v9Jzrb8lVGjxUcNwuZWMJc4OeKbS8BlCn7w2V96el35fJnWf+eBZ9wQ0
3V3ObO5DlyAbsJxfNY6C/VOCmR/IRX1KnILdkBpM8qqbbFTNMzXTEMMXCr9T7aod3Nw1wjmpKPv4
DFa9HAl9pkMyhBooFm4EfkXDxG7qBVKEJJDOnZdr9O65uvLf4EG1ettoUMax5x1mrte3HS54zn+p
p1EqAJebmrTUvvnaI4vRxT0ifspLktqLk3TCvRez6YrrgBzslupBA29JXRRS4UWQOTRUoJqIVDbW
7/z3POH8LIsgWXGnege4hvBA8FcjLu7DuPx4CW8oAL7TSm4MCfcZV4KlGa+DaF0IyUVpwNw8Bm/R
aZWst5ifbgs0pBfnatM8Pljr8uYZzpuOGVN/O3eO/QcM1ZY7zH+ApVXwt7cPuLOrjOlYObFmbWor
ryuWZYYJKX8HSKn2iJ1XrrP2ZwW9F0umx3vKlm9OeP/gVNHPGQbTWNm1YcrKgfXbgHlKW+82vRiu
geTjvy5M56Wk+fjvIim95YzsyPzxVRKN9KcwkRskHwPZ4y8xBpTQFUOyEYgJk5zuMJuMUF1DAVnH
iCP6ytJacxEGhf69DHPdd0oC3S8AY0fK55nykn8bibrUbrgHEj1tadyvL9OPaWaObSAYDpFFBMQM
faLL40a0wd73Tv4v4LVwxhPVoIzqL+/cAOhvu9LE8yb3nrVPADD8iX9TmDNT7nFISNtRZv9au8L3
ta7XkqqkAqGEPx1vHPaZ4xfx5rJZWWujQ0xafuRcFsvmtyo4JporyK3pD4IuTol/dHVzfMMzgTBl
QQJNwLN1s2qLnqMzlSGK8E3tfchqo7M+hKHPjM5NUuuF/Ec0n/ERjT2ImXn0fgJMIWvA5sU1Hsa3
R+lw2va82lOYTv46DkPPpcXkkWYDtGPYJDhtD1yGf83ly2Xh6FcS3786KBpve6j0giTCN8nboBVV
oC6E3OH2shzi1kTyxYGwSVy30hPJh1AjZPDZskabPc44oohB1Ic+HyoA5t+05aGn020S27aHFMhv
hJh9rtEB+vpZjU40IAaQWzaiYYYgR/+8U5Z0JGUtX8noDhvouvu6TWuAtv0c0rNUfnsnBkBYahY3
Is8gKJdiGcXvbxG/E8BQXRiprTVhoKpfihOkzxGOP4xzlkNkHsGnLYyOvIN6PL8hi6U8F+Vq5dvZ
Z5iwqrhp3SjNv+vxuQQBXEhz+CZu9oIelYs+9vkNH6qS0LPcrJf0lrlQbFkbDHeLly2pYIOOvy5+
40Sv4WZYDtRaRdaR2yo6yiEgaOzjM+7wPey843HoPhxDcRAKWcFqt5VV7E091y35mps4LcAH+vrH
Yojbmdsp3IewG8q25gZMj9zPCSzMaMVwWUbTwNpujztqRGHJwV3GlOXtr0hZdjsmIvt1I6bB8YLs
xkd9O0o4wsNd6HwTzxPyktGHeijRxzB+vC55TUwdwrNC/gVoMDEkIpjFPKi+3PBl9azXWxwezV61
mbk93BWGLgtRTgPNhf3XgapaGPldN6QC9w/zPNPGjsCWCZZ/bYgQUkpYIri5vBzzOmdMpU6OXdZl
kpWKOd7Cm0fppMcXNgOakAmskITCXfvsb1/nqdlvbZsh/FCZsb8V4wkSlRad/CD8dkQ7VrNyWL3i
oVZLw0kOwpt+TdRE2gaLaQfHpfC8xdlj1DtKhNzFpdmjT99/N0EHIsbPf40glZm95TUG4jxUYxqo
qh8ln9BIZyfcWw3NZClTsN+LLqAkR99wIRZL7JwBJfeU2UzP8yn9j9p7NEjgU36DQQddzKJfgLYk
Jk1V4FK7UX4w2XS7OL3/XPRZXfDZOMOxv1S8Tj3CrgWtdkEyBJ2G++fqtATQGh/YDzL5up1j9IuF
wilf2rOzwtIm/ZrKiIJv4pfq+HGU0X6/cmrvL8C41PfyTSRJTYpZsxHRfkXxeO/m4q0J3n49nWx4
98/uQjF1SE6NtyScKCwVHp0k+XhkhZnESYJxlLRrJL3yEn19c3O4WCKhrvzithhrQ9ctrZhrELnd
8xDZBNa8OlHzr7U43o3ZMXKWCEoXCM7/gzrlyb2n/L1wYgNrernvdcaE8p8BIdtG34lW6bxhtqwv
WoQk2oVNrad0/41SongmWukqziFrdc92t1bT4fU7ETe/uudQ6GvlcaG8MZlOF1cZyYDsm4BIY75t
2Jib1mPt5CFKdZlPQqjOeqUeIvxpd5vvLxpoQUPopZRZLTsp6cSHu5gfnC3UQMF+6SB8UV3TQsJe
auo/CBMJXHPUIJwpFNLudxEPYTqJ77qtNlA2qAh+0LyhWi50VBPbmP6SHfjC0uUMGadNr2WgIboi
Sv4m7PXST3P3PpGitp8ozpeQbjzgh1GGmAj7PPIcc4X95cCSltnEzSp63i8TI+UDzhFXKyonfKVQ
Bcz5f6Orm4CUTB4T/Z3szDtgdFOaQo6fAe5wuoq+ZUxNSYvdSv0jCzGy7ZTKQgcZ/5x3E4IhcZk/
1KJ0EHJg2z0eqMJpuxAwlDjP/c4BfRrA6JrAYnJ+Sgj79FYH0FEVHQHzRn6sTpIKi26kC4xyuIdI
JGa3RZWjexWJ9W4W08nd3HugBTj0PogY7pePnijP1QEaOEhpyeVp7Dblow5s7q8e63JLNmsPgOV6
IRr6IJnnyOBqrx5n+1jLb59Wua6qql7uV5d5eNmmlj/dvCgsO0ZbAzWBma6VCyPM1QmOuM3dzERO
2506zbGs2hv47rj2FtYboAmM7Q+5WayoieiuBk0VG5y7YaIdsmJ/XUXjlud5xAOjYOkeUdZOAseE
PJLaIMkl4rxnXw+9LDTKTzt4un0/zjjpzWNcYIy4Zo/lN+2nrPmBMPD4b8P6dsbb/Pn2/TYJF6Tj
M+4IKRK4QTz7EyxPojmzM7cbs0wKzPGVTBCZatFYjY9Ia557faz8aAPyndGW96aXap0KEumjsjyb
ccdE8I2o/HYoxbi3zMrUSCXSVb0f50eUd/+4l+Pife363JTmEy3jy2sXiZZa4+kozZS0CgbCEq0g
ZKfcPojsOx3c8wX1/c/YsH1lO3jLyfPKFbPhGrKBnCx2e1f4o7k/K74gz93tAeopDpsQiywZ4dNr
64gZDiIqkvgZHq77ZtcqW5tXgbd0e+axUo4j5ybvKDZxytf1zNKj1BjWMHxaIpr8R5ah8nJauEP/
QEFgVkz00kLhst7ysWBiWyQFcEuo6H4rw842KYPiRori7Uuv9yyABNoOiFovfDYt/vUtjica0eoa
QxkEU37Db96LoDEk+Z2nQ9XygnPR9gl5UOKUhYO2QFpSjI+4Ieoq4QhNtNI2RvHAz/UWd34alzr3
Sm/ljVh36k6s5tGniUJ9SSmZSN2u9NXShvcCM2++vVamaEvuVi+52Y1BMWxwcfIqzv38OzbwDgia
eUzhr6yHsa/NEB/HWRA4fBa/mOlTCJTt7VvgoM7Gp9hgRoPq1hq7ZxP2HkRBFIFGkKQbRRE1S+o9
Il9AEtypL1WcUQTlpRaoZJD3BC+MSiywpzep7Qn0SEVWEY03ICyMFkOIS15H09zAHUjj9TbF9fwy
TOxBldFvvdgUc7qnp9rCr/egv693fuEkifg4FbF5WPUuu9ab8KGCmuf6FWmbgnbzcJ0IEXKqo8G2
s8tOVrzNIEt5nG6GQiaWCI2A4SNxUHPvwvCFamOtnExElq7EpwOSRGK6bqM7qBRWQBq+CSZMM7NW
GHmv/U3RXnB5Xna+JjGdr50IVc5uZ1HpTYcReGt2rBMO35wwrtW74OVmecBvHvZ68K/pC2giO4fM
XE68xWZggM5xdYtOFlHkmuzeQGfnBfoKhA4MF7gPrQr1NFnCaIPCMphrx3qtCrPGoKjuCYVrDXsa
GTCKL8qv/EtvM7AO894HCfERwjnijANtRY9p1L3wGNhWkkMViFnCWGwos66/GbT6pWsnHq6bEKjc
ZxY/LLpf+1xvgW1j2z92nTclzbNrQHFxIO9El2gRJ/Bq0+S4z8CTmoAButkNMQxkDvgh7/ijtF91
6R0QFG/1OjXWbwXBYzjbjpuh903peWRP+WTaVOerPE3ITjhWzdEfzWrky5tNs/oQQjRYi+GG7gEg
b/xSDUO3UXXYJ0GPTs7XksLRxhYfILgGhzQKaurQ1FVOeP8CxCTZfjDbQXj0lhT72Iilkt4h8ykC
dZIdM64kVppGYKjuulwhzuN29ffOuc5FIVHx4SnhveH5fNynf8YDA85Jv0WWh4Y5uIWjKyASbQdM
pgv0yMLn23Eh/QlSAyjAAR/dVlXicFg2ZRbmMIc0TVy87FuYJ4/z4tqWP1zPGm33M17lFUN7Fkr8
tqwe7SZ35xRaekYMpiH/VJE+3x/JPOKYMLe0j3jNOrKtW9aTBI3hcNgR2hg9pZkjaSWAV5m6u6Zh
q+SV84JnUh9m4ccIp+n0znaPX+4O2QZZHBlSm60KHBZzjzBwn7lAgDBlhyAtlzFZZDv0owsZ5ehJ
GjDdjkx3Rp0SzuRPAuxvo2ZJIv1U7zz9OLc+gyg3okczQDV63FJYfKL9CFCtn7vEwjbD1ca49adZ
HTCb2wVA06w5TTUu8wC8o0UXQnVsnBV8z3BnIpz+r+lQSTDWhNBXBsh7CR8tsXVpFbXvWEPcqgcU
83vJoYLx6iX+k0YmcANxEOdCqnMzetRLoWq7mLAHHJdZzgpzivMqWBPuk5S2WOJGpUJmwDYfdqIO
uNWI9otymTE2Y0QeGXlwaiKqLLFf+PsKJFtW9M6SBHtC7lu7nODGO3YkBwsUqu1rpqvi74/jzFe9
YiPofJJLnhUam2sm6morsRgj+hL+5lnttDH7o/590v9nrZPNmS+VeTxX+Y4kn9ngFqMtTubUHXxi
ZM+T2lR21MAQ+UbpTtpmJoRxnEjlR8UQhnqmgSNazEAw/YluRDnniVF7+8cU4TMknA74yG/Q03If
XId9PW/wQWvVS3mZfHQOE9JHDD0LRhK4sa6bOVEjFD5Jumh5oZ/jyY9HZMKdTmcwyc7oFfsAng2A
PkfkY6z46K06DOhzbBap1vI+w9yHbTGbIMIkUNx6YyOjg8M/+BoZKxdkUtVpCcACZz7nh36fZYRi
i/ZYWHUiJz4dRgz6Hpc/sXmVkpI4c1OlwxG3OE2pohITLAmhtVJ/A/GmZJF1J1kP0uyzzoH9n4po
Yen2XMkiDIALR959LPLhe2hk+u7VqwVuVMSeRzSHBPtnl829wJ+1IcYyzh9FLvdQJ89J2FkxLPf1
U8nrkDaPo7VHDt2xg0rLgWsZNXtb4/zOnM9LDh5mdqGdZeahZFmiIMVwNxa/AEf4D9XwvYv8eIWo
BnlX6qgdWkQNC104Nk2/TU9TAF4cxiR7XdUrT245Jgs/Vt8dNhpLjHRmvevDkcWIllIi4tIq4YmW
lXiwDAEoRK03oM6h9jUV77+UbZLsrW2i0xOEWiY7705fT2FqA8owEaEWM6Fqjmc/CX4gwyOkdksX
zvpJFOCGvJyK9qPxp5ugs5BLBD7ZxuMm3n56uqBToexVL9USGe9RH9Z1ZZkSxEGALacbhpMXzdA0
xnIaiqnDC9a5eAQ+3jusIJg0Ilvb3gzZzNc7WvzBg/Q8+vomL6tSgsfb0XAAkdoy61eclMc3iT7f
fS1Qds+0t85cPxGH5vIgi/mBEmoAg9gNPhlgbrCg/HeuoTRPQEvIuUP/XpSkmwSQuUIXplhjrsRU
XFE/39nzz0LwSSHknvAutP+XWSnhzxbx9ZnAoHMtKFB2D0bIMiiGPbfBQQhCeqtHUxxYGo++qvD1
1UFxz9ESr5xYalXCL9iZ42Uf0EhT5i/nw629LPa+Jp8PsD/exUVyhLKFqizL/mQlH+PGKiXwUDal
+B7fP/ZUwb3yXd0NvGOsPP0Cu2Bsv+hTe47h59//vWdfreHZvcwvF9dUnP7APdhBtdFj00hwExEU
0R25M33vESh0QrsU50jYHQesrzKjo6FiPCCYMJEBYVHobPM+DdumELHiGrmEO4X4F8whQcQGWsU0
H5kgoaZYgQlqdvP8DKVGR2/7eY5UUrVH8u1gK5jU6y0FPGPwOnkaPe+/T5Wagsw8jt4kPQjocjEb
KZ8EIBycckYDNELUuDZaa+yzVXj8uypBjWkfq9mEemvxJLm/lghp1nE7tttCaYUfAq6piVWiidcX
eo8rO3dC08Y9xPRXFGRZhwKR3CRSybuBoVkKvaKBmm5LEYHv7ChBhxU8J9MxeVVw7a6C8FFCAkEu
siAdBvAuLDia53k47J6O6g4+980QKF48d7RQiHBYyMa0s076BrCHo06C+kCZ3QxusFz6a9ofJeeJ
xsxUjXT95yrd2ZUJaD24jzADRyHd8IIF3bbiq0EjOHeFpxnD/SVIegS4hFB0pFNiuHMe9x+nqDrc
ct9XhjgjEiN+6hJd18fbWXSz0LZ8ktvoytnNiyiqXnQv4TM1JMyjxk8gIQ6qWUdB+RJ/+S4HuaNP
o08MjZYlioM9w7rx7dNlamO6letb3yonIuOVSxni6VC2uSshH+NgFnhvhTPXpnHARpg4aDkixLAb
wySksQtpzxUqtgXxXh8E8Dd1OO4fJguF9JA35YLU9OFQPOR0aRf7w6ujl9gKdTGyWVzraFRAowcM
E1QnVwsN/oCl212JSc6nesHHFxBNV4/Quc1GM89qahUGMDTx1yFSB6xjQs1ZN75O8jYHG9DR3DPU
qMWv6UeJLZj1TeqD36ECMAzGxR+hfiS6JVtGkVLC5zMy/IJ2HzAKGZIdI0WcaQKtt0T5E0NLlFxA
muuPU9AY9eXGO1j+9z6atGZfZLRMCWL4/BD1Y8DsLaQIZAe4yJ/gr4sYl2q7tcFodCkTKcINHZgp
QOpp7mOx3DBsB7P1F0wC7HZiqJw3do+si/2+AfHhGtQCozHtLkKL5hf5ApXiF3JTmoSORF+EZCWK
j8w0hqnAFV08T/F8xtiF5mRkNeshCuEbyljMTg3J5fpP1asgnEIpGUj5cxYpRZApcYOvNAXRC7C0
MhVp5qNmgzr8/2Jgp/o+bCqIpZwlRxB8y38PkhpGBJ4txhhrTHcrBd6cTRDuOhiDrkdu5VJvPqar
bdl4GDy5N7oG+cECsG/rvaIi7CC+f0S+UD7X8eA88rmGDBoMj6y6hjhu4JhWC8QAIBsNhdBQ2sS6
nk3o0EKv/6pND8gM1IVFVOgVIlSDrOY8/t7S6cE/f8O4o+IuYZBKk0gsatSc9JhItVSxkjc31paH
588YRwwekFJEa6EBFr8+H00dpviyhpH1LfSK2tLdXNMNxS53rXjwKfePv2Fq/Lb66nw1Ry9dMDUE
MSZxIvsPhsX1RSC4DPKociLiHAPaL10QOhVVLSdLewGCxAdL3pSYpc87k9/fi15YqMvv6iF0bJlI
yJk7wDezC+kdcFa0XFem3FzM3zi3e2R6NkQIuMjQWo6T7HhH8GfPA2z57Vl7NfmFvrbolCp2BZWl
HbzRnubGs3rwq8+CrEUYH4yP5aZ/ohjHf/I5udxDmIJzj0tPXK4wupP0D5FXxfVQ0+eIA0EUP0dG
BGIm4LrK5C7gDvBs+5q7Inkhf3TmQgzrifaf02J3LBA6V41KOlp87eWzfFtHuhu1x/VXQEKrDp7W
GWLZPwlEc0AeAYTdkNo6So84yK+qFI56bPUnwFUGhpaV2ExmSucoC8JZS76JDtUjGw7t0kZydlXT
Ue5jTuDTd5QdTGzl+3wxqJptQRRjhjDrw/RxlhA8WQqhJMUKZEy7TPOM+Irj40OGerg5mwHZ58EF
d11hpSxhfEuluNFgyfSC5yIAZrBhwipx9ZwCgn2qndwHDoNWHdC5einoRD6FE80fp6QOXqlmI7wW
IcQc8GlDWNJJ6D7GUn63xOtCxg57/75hxP/BVYltL3IfH1JyIWByzQ1OoeRyzcS/078F1nB4PwqP
mEhw6viTxLoL6cFSk7FBxhA4csTbdTykivwqTxzHg5bPS6Ag3Cp6di9VQ+zpU4urXaiFESpbEmWx
XpNWyaKVcTxjPnHoQRDPK/ie08USBiPxN2dIIdEGj1koIqnVMZpgYDf5dFF/CFg57LvBWR2MZ8WR
mMajWoaqGBtGcJ2owKeKuSyrSj4cJIdIGHlfnHx2ZxY6YFwuaAOcwVhTpJjKD9DyLTOnvFCLQClD
6hbjpaP2iP98hSIYAZGmu2707qjcoe24pyI6N7o/6jm/zVqhaWux5Y0SGaPMgjRivuxUe6WZznVT
2IyIKMrkPOYRQWiokYTK0gp7+b0XjtSiiMsO4IJTgeBIls3h5J9/c46cA6ZXQ8zFsQ1A5zOCEDCL
f8R5lpmycw+bJCktiUSxDgBWmWwk6a1enErfuhDmy/2ni4z2QhjRmj/JK7HQFAati3JYtVqCoTHW
AvqFCx/4OxfOnD7oNSSdgA7SQ9H4qrXYMq/sE93wuiDmPemN8tFUDuSFE9aEHltehp0q4/B3SRTO
zfIyQ3+zz3CvjbjUGqeTrZSBEgNK7Zb6xU+Vrr9anwXFZoIYBGfbh/nIdMcgo5QSpUk4gf9pIKI3
fHXYY9C9kwq12ompxBcH8e3OljGHy8qrfv/OK+barXF2PfJlsb8LF1Sl+jvq5YJCGpzyYdNFgtOZ
8J2Njsx232smRQqu5iy0xQg/bG0lB0KEo8YfFYW9bcq+2iOu6Mm787UvOMZw3ujZN2Gj1zhfr6NS
mHRf9/8/piY2a4xxDpGEBcovUxolzQnOHyNvDC1g6uyt+z7yjZoDkUF0DmKTWJb1UdWuTwdkqlAn
ky4Z2cKTe9bCAok6F8MCt+ylsJQuTx+H0Q8nVQZF5iHe5OAZpy8Go72OhZ/jvz7sLMrWfvg/elyZ
ZLBSZlQevBDPtSe+pgrp2020fbxumKXeQ1L6iCgytb6EXiTQTPRDM8xQcwQOFjOfZorXzkvCACjb
qcdoHV9GTfVsCUeu2VnZryKR16FmbCZVy165gayfsNUa2pDuieoODLXxmHHn1hmEU7gxJWYaDnXp
9g6BO5XGXejDR9cpl8dpNKr1iZGLOBFJFbPVG+UKxBMgNFpO9PdnTqcNCJ9wdCC65yAU0/FzYwT3
cINGRnkSoBI7CX/a+WtzVGPOSuT0LFBkMXcXXBG7LcpsZWFJB8sHELMeyqxPLh9msHNN/mR1Jn8N
Z0QNrBm1wYuSeHJuBbNw4cBpM3xEy51usC/llHMbzxnnRZ7WWOn7DRnQmdWFgr/DIbcwN7D1/9iH
bzlar4oEqtg0Hfq38Sgvbr9EoYKItUxCo1/MamtIxt7GK4tjck+CN1K7A9UiYIebgKT/P7WX9AJw
6iJ0mZ+lTsK65V8H5iPIrjUZ2NCw7Vm0mudZ5yeSgS1FWajQ7mgPiQwULl+H4uZRhAIKC/lN3KeK
nKNR4rTUgju53pcF7WeWP1amRtz5FRIc9ZcuHSdVJPCqCgnybPsMgJHZ6wf4vosy5rVjN3CIlEdO
KSprj76VMK3JpdMrDX72RidgwVDlWrzrTPp2HugAqKQ3yTW12bA/IfAzQCVEnhAsiFhRQ6QbaHEj
w0pgTbxsXZej4CbPWaJwv2JmOMZPyifgWc/jHscOoakowMKOPvxaHIsss1IaDrsr1bOrZXEYpCIS
HyknyWgS+3IfMYR0xkHd31k3gxyD2mnyahwHhZEc896zFlphf3o7VzK1I/HDL2hVEYlzwGSI7HO/
dwCR7wJeyrUgiWBOjBWXDTAsgOLCPySqaeBEOpBwAhv0+n3GkQwV85lYZkm0HCA3c00cq+JR/Rmc
3UOHvxWHIM1TKoLOSwvndmX4OUuL08YIFcFNLmnRxwRf3KAxdkYXeqESafhsja4+R/TI+TTFJ8bF
arNYmg1GzHmZQqhWB+uWKmk0C1Li6JB2SzSZnF6mRFPgXuoz+R8c3kpUddF5r0D70gno7OtJOYSS
rRSb5EGu9BjOpzoUA2t9qPlvaorHb+P/qdalFW+KkA6Zsjsu0ITqNOL4NMClhxuotjMzOtKFZ17j
QMevFzqmvW7ygdleGW/JPDTEXfjAZt++6qqpF/9+ZXxhlX5O+zw6aszFYr02bcGfYwxzMYgXlooi
cF1Pp5wiVw2/oY+pVs0GOh6VK94QnLMlz4u71ZIfktH5DBRiSZlSndr1dZDhJ8jXNI1YwNneE5QH
zqtyzVGXRtkH5g0TYxQYeMSqvIsA83yyt2VWkDTt0UFC9xg/3RFs+5Ymzq4BQy7cxMwTgLfC8Feo
P59AYzgmwbKR6x/nMRljHlHw+BfZ+AuvosJq9WqXie1cW4Kx2I9V/jRRZrPIqZVnh9BUT+ENQkrc
BU4ZYiT54eXMPij4C7JhUZxYEfHlkQJmgfD43yQzl2ejmtksRh0JIgPm9fCBVNtPc/9y88rn91Qq
ialO8Sbh9nt/LuaJN/nXoK2egpjN/W6yQwe1L9fXCpI4YM/RoXGpx4yU0PRtXwY7BvltX3cpQ6GP
XvTcrdMbMYfoVPVf1xtbw2EUAYoxOMqtyUtVTJ+zCPJ9WRe9f7FYtIPy4afDzOL1+3hQM54wiqyY
cp4JOh4zf4bcxSkFufp9GMyAOXkbsXqc0BSFnxkAkF1rrTvlsWZ4KVoWrnzAUbjWS0rt5NvkEKny
ncTsjS1uqHYrGONle1sqEycY5zypTcKET4Z6ifkVzeR7TQufyqzJC3dgdnUZvlFI7ERhth4J+GEQ
sJSKmY+Tm+wNXwGFnbe9h8GBTC+U4NaZuptKbBnY4yBrGOhFAE5oZqQm9XyLThqRhA5POur2NHho
GYZ8l1i7ZjUUMqHWUJLGepIccF52kxrnRVc8gQmTGtkvk7C3U1OcWLRJKmSskXtuQHDcThYEA+kW
gZSRADpsJ5fssdHFV31fHZ/HgqRduS8SBz59tBOgdZlc86jsHEgajEPrCSmGoo8mYNNLgwCFrOzr
JDpe/MV7V24QaZXTQfJXlXn1fh51F6SsJ06fHI3RGhlbb7ta3yJe5n7bhxDtfD34iCRuZ90cdgXz
atsforn5vcaWlHho+/d0jTMJ6URBm7EnLpOR+/DbSlFbR97pjAFE/r/HzI8pCok02TJxWgDTXwHM
2EpUs8mnqxIy1ouDnB3i+HoIlRpo+Z82ak4Foy9FQESJp5JDWSqeMM7tUfmKPK7lBvmacNA+Prir
3Dt7tJnFxGdUQ+Q7VAqqngS+07/g3SRj6RBWwkX5ic0dSJbpe/QbhWbqwCy9FYrw/m/UcVWLu9rc
rWxmHIA4Ru1UkV3Zh9tIWllC9o04f14SwkySNTG5xDydAXELuGzdNEF/fYZPhKkCzcRZ3Zeo3Ep+
NZ+j3PzHrvMyARUzDfEYqD4+J+tN5Wt9M3nbbjP/R5nOOcPllNukOKYm97N6X2T+wZZoi1F9Zn+k
VWnVTx158DeD92bPyR2yDgTq0gtqMqRBQfVUMjOC1tu8w1/rnw75j1MzRF+NcZnpMCcwH2AJNHUR
CQUowfSuY8Jgw5mf4CQSFwhznY5bKaVpxgK6A3UkSHfcAsAtQqaK0vNuyAh8qKz8PjrmRciVsoxk
M1ptlb2y7Eb63zq226kYphcon61bE7eCHOCM6SvYZyTMJsxa4fzJZwEZUZ36g1JZVREyoLnNP9qa
MyEpkPJ6mNhQIGBkVWky/XbrLm+sfNi95zC7wlOT/7N51/sT37xcnYuIcn4I5CevpoatzoMxBqUd
vOJoM4U8zgWBZ5s7cbsoK1rVIUD1EJyTFaeeSZ9niZY/rEzi+Jd/eatwaN+dX3W1vBPpZAusyBEO
zASfatXwmjBpNdvRN1mrDLnwSsG8TzXSrNNu4c4vnp7Q4BQaFCZzF+dZdPoe7GquWZJvTYf4f+Y7
pLRKj5nLUVRyNIl6ewefogURTSf5rKurzV3epzChDoXRXYjpiRs+pnOqSG4Na2n5txNn1HEe7yDW
ewIFtB815HxU65zjIS/hBEfMFA1bwjN1iC9OzSE0aTx4NQ98IDto3EEHFvJQrq7P7jsCW0ej0N3k
DAHUTfzhD6a9lklu3RRAMFeFnsmiaxj4wgT3ew/q1m2Oo56KQIjnx4NefNAI5KgPyd6KX4XgiRIl
lrlmweqYjZvLrAV4aDUPzbLrtdpvWkLBR+4Ut+5iD3Q1Z49p+k9nQ/TzSCdojSO9ZhFHYD9lE16X
Mj+R2UnqQbNdlGx/8lcnumqYmSAWLEQkg8GFnWzL7hpakvbaaZNTuC/i5wa6PqpXZWUGwCA7qgjb
Kbb9c0Zz5xXQJ8GDyo92Y+JaYkti76WQnfe84fwmxvLx1fYERD3meCptAMH6t7mnLu4t0n8vL4y2
1yI6f6geo3K08WyiwaBzzOXvOk22c+tmN9qteAeBqeOqQX+RnZfDMqoIJqwXYxzYuXNq6eoasP5B
Bncx0xKs6eraZWaOzdhdzRGItW6xPmkLEIDdUZ6dXDnmDWpLtwnajkH+Q4dPWNM8tCEX+wzBSIkq
CZV8WNVfJ4gRle6BiLsKO2u+MzRJI7GCDBalM1RqPHpHV7JyZm4GpdlAmYNhnGmCvjVq0tPXGLRz
hQ7la3tnFsGCmNuABnYKx8gwrfRhYvrI7V214wJl0G9rAhonQrPUdlCLxqRuo+e+NFDoeNq46Y8/
AscxC6/xEXd0x3qc24cki9Tk9DEcx8LitHOshmHHGT2IbsH0EcR1IfmtuCrYtfBhLJYT0lfoornD
5tOuFaxs7VsDqkodj7dYkRByRRRB0+dJvkawcwrI0qHqFH7Bs46TiQObHVNUCzuhLdvWHag+Suve
4mQATqR0/0TO48RL8WCCb/kBFbmwkLL4nIk2tyJhjinMqkz5o7vqNhI3fBSZAuzAhvkcTameMBvE
4guXLBZZ7KWQfjV+64kUKXyHnN5FgJNKzLC2zkpv/iukyXEvrjFHX65vej3e8knsAlZtStZuMS6z
u1y3NeRgqYmQ1Z9uXSjRpr2AuPO5iM8ilUUd9/D4wv//kW2hcctymxoKP4DfDnSunNe4dha6Q3Ni
5K/yxjj/h4N73cmTZz0HD3bM5/i5YM7aH56SHFQCYSgohAytQ691lXpE2P8lPYdPtvNrkPOWFLS7
n66Ule8O+UicfF2RJqxb3O1NZiRSGzRwVBvnv/gxEzYql2lDDzG6gIlkSf10uwoBSkhE/OjGygYD
QeTSBviImRuZAa3CEYmEd9O0lB3WNRi1W8Ct2a3arlFtq98ZsNjcDsniDxUCE6jqmXyK2F3Lxv1D
CTR+Ya05oRYi4XfsuQNXUTXB5o9cQuLfa9SFS1qgqTvDWUw4YRhbHimM3DneKNCKz6ide1WRe3hM
Rx16ClL+FbW0s1T0UD5HfzSaUxX3Qo6CeBWU2vp5K/gflDWSJNVkukFWcP6cZF6Ei+19oxCb6Zvo
xVTXyRSFOPrJsN1+eDoaZqg9Z9U22tuB/kNGfIGB5TmDasUieQaQ5mPpsjtG0xjXOxV7bHJ9QJhM
5HTmDAhT8aRa2YkDZHOJ50OeRgt6ZNRmVHP8fG3h8dTSuCks9uGGpXSLgLcGa2aFFOMWXAVIaQIk
ASGpZcO1OPKVEEjw/cF8hQkRQJgnYnBiNTyo0lMWf9nk2gGJv+KMcyA7GaMQyMa1Uus8xS9dqCGB
mXg4z/SwZTy+0mvLeTPT402d+0fTI4zyzYZ2OQFr20Gp1e5iStR0902DARGJTNGpfeCocIbAZuVq
mf5TApZCFAULOsmcgmWiMZ8e2iuFlMUZGd8/6xO88jH9opOjmZIAvqr1QKtZ6LqpkL1ldUALzaI4
tnvlunYY/t51ZmtE67l5cpqhxu3vf/SI8iahAD8o6uv7YBJEHZG4ss3O8GkcCmcDGqjznY/3AP2U
cgtD0mKlIWsS8jY2k79Bl912q7vEXgOwh+shXP6rLTb7ef8xZp7eWVMAlup/ncnNApmqNqp0jKfz
1A3PEb6NRxhTBnKAYvWwkxNiD5jNGbbHfzyYcTTxgiQTydO3Zfl0QgjMvdoJ13bY0GRmIgpLTPqx
+l+wCdkqkkcH3kmGu+yClQPCxeuL3PnkZUMf2E787AW1XCqf9lbpD/cEz3kATRpTzSpN15i1oz7L
j5jtZgfBG8V6jxO3X53XfTD6QlnFetsx9hp7HK3H7UPa7S0pael1ObOIbBAL5UVlCh2SK+M06MRl
MSzownch1EvCVMsCCkJXYkF9JUaVjFHhzl1w+cUVYKXRSNiuezI/xbhv/d4nnxURvoyxb6NBfuzO
PJGiOiCCVg2ORGHW+FtkjRb6xw0qQTsc4GFq6z94hxLL2WqyGV3SD+m7sWNLmE9YaWg+eFqM/m6Z
nCPxH2QMT8ljoPaeewFsZFQHfBWyC9nwrlhsGZ+qDlz2MSdBPwmnzecaI1RcYmbryGnqsgh4tvy2
c4IAvKzlRhtklmDu4HE4s7c/WTG87AedgMVVic2NwAfCy3fXZPULjtQe6sflmdAFVZP2Laq01YsL
VUY4TfCGnCqr8LQEGRSB2JKFiTdbmBPDwInlEs/mFw9dLg8DqSbrbYOIX3kN4fFv8qebTtMg/+hL
u5R6Xte2qWcWMbuZSYJzzSkvMnCeWSCi0wPz8+BsKI0cRBrxJqAjpxb67MD9d2JkHk8NO12ZwZZT
zOyapdGplKt3KoyMEsUpI/pDPW1nXLeo6e9ZGeJZiKjoN9GWrGxP49mfmZLznH4Ha1/ScUGayHhK
1xXGtQ62TtC5gNBMUctzsRkid7UFViDDPRKig2Om+hOpLFTSYkNU5iRjqUX/Rpa+3bwAxryLi1go
2rJuk97qJdbPKfLA8W+vv3e6xcrHagDuWS44A56EojWhpZyqn2Ke7ZFkoYQmhXUM1pKGKQ7cxMWE
QrIGS1yqPJnXRQ9tiLo9QnrgWsmjo4Qf2b6aJF6vsbUaLGzlZUTViliLPTzdsBl0r94bbq5ECRiP
wadc/trEjHYxpm8pqskuXlDgszHpAUHM4LXsQnCt3xGb8yhvBfwfLFmZlBzv2F2prQwj+zpd9scV
JGgv1n5XxrCfvlBbukS54oEV2yAE5L7HIFvbA2w+XYq5d4EAOSd3s+SjnvI8tiQmvlyxXMIPA2Sz
E/5TSCw9SG63grP30LkXs5CIgfGFvaoJfTQvT4kdj5lHgSGErf6cIbuvkx1BeOPe+DjsyeeBDxb0
n3C9i75T3lub6HECJfwz7lAkGm2hJ19GGLAWHtpch22ohBA7aDKYjV/aJtB+0qBhQiefMCDjN7Uy
opHaTRZ1vmn+R+nlfvNP1/I492L4A/QsHNJONar+Rj1yMhHaYG2CNa4mp/PDQUH/Q3z0+Bvwjwce
dZCN0YW9xfa+s48ObpAqh242H/SK4j5Aj5mIpEAjtnnbpjwnvlAX48F2CGUXklo3Rf6fLXBYS7l7
fVcbwXnGOiYxdqbgc+Idlx2MUNie2wXcfb7FysRLheEc+oSNvowmqY2gzWEWWUE8MvpZnUr7qnVS
R01SurKp4o4fel09IKg4DGGp1RsuEr+KlZw0y7R3UPCj+MUioaGA7bKsgs85+XDVvPcbtAGeTDl/
cYPjhQqwJYBB6o0P2ygpymcmqNb2kJ/FX9Q5IUFEnaAqD2EjWXtKs8pK1gs8VQxSaMV9jJPe9sJk
VwMul8GWGZGzdhzV8OXSgBAqT3LlKskY/RgzTEmnsmLVnizr9/xgkuPeOhqvTOvKFqZ71eLv/VFY
neQO53JNKrjs8PnHF2lsesTTlkdGc8lXkIGvydZn3GFwQMwXb9og2vqW7KWN7yXo6wvmtS/tdX82
vkyx2i9f6AXdGFe6BBKyK3cvUEAXBDA5kA1vI2dgD0I3fTKBiQ5yetS7ka/CNEiLpbGxsOwTky2l
Uknfzo2tTDklZ3B+U4njiIiX+0t6Utg1IJbnQvlV4E8qOPtq1pnffUzsBFe0Rgphha3QV+5CRBqA
nmDfjcZge9EBLb2FQMETQ3DGoEiv207Xrsm2UsA/n3c2k0fiDxUzvkOVJNeVUCMmmq2pwPDCfQYa
4gj5N41nqIEsDblt+zMvG5WAXfoc7a3wUeFUtVH8prYJjyPrYIrWKSnCVgpCZGVE3HlScdH3OeF5
DcdemAq1iwEBd2Dp/Ya5vxjm7CBA2Fg0CshLivCdP5angne2vU695PdKTHCDCygta0KMkCgiyd40
OULB8dmLCaNeZNi/TQJGRNNE/e3+sERZ/gI9zCARCC/iCMrDeOt0y6AhLun4quLOMfZ9QiU4f2bM
5x6mLka64yPPXgv0G6kXmFkf5pMRqCVKfIZ3i/tKyZKuGwTP+lYKmls2ENThOnJMUaRE9XLPoyTb
hu9HcVfdRxK4Tkh5/aRWELGWVn/atUnTkylFLt+68+STSvfknzVtoNATOqwXJFHEL3bim/WT33AF
9rVC041p0LaNfztt6SYlmipatFVg44rMLLZKsBA1eRjQ9Qj2UBJK+Bjo0PSB1lvSCPY/TtVbU4qF
K57ec2DiEHBkT84i2JkvUrj5yT8mVUOrJpE+9RT+AsW5eMAMrK6JmKEXCHIgJU1a1943bp1Gvr+c
XJjA3WcILYzW0Soj+7mTvPiYcOQlFlpufec3VjBA5pwmP8nH5M/f83ZuOcP+iG6abJ/Yv8x5+pCk
ERZStei8vt6LHCsFy+YCoEd2frQjurc5J4za201MrilE+g2+8khHn7/vuYSJX7m7Lm3zP/Xf9Cs9
VRuWDU16aY+T8+pCJx8eDWN5ELx6lth4P2Jf9Y6qr0hS7gRca1jqIU6eDWpX6o3QqFFAxid/RGpK
NGmeYkmzJsX2orv5zT4+Lm55VyKOYEhlgQt+nSlFGQxe6DdndB7BNOgafUSJVzrmMOk07H4NX8zp
GLlb/LfJXZoaX/DmNwmFPJp4lDIXqwwpVozdmENQ95OkLLvu3QkfDQobFs6RRaMDq406X6Z/x2dd
5b8dKfzZeGlgp+wCGddc2LHsKgV/6eb5dtkvKbtWJQp2S88g1n38G+9WmSA/gnY1pX7qOCKE3RDs
DF3Ir+x2I5NvTeFAazyUuThZ38ECCogCVrF4aqv+Mi1FQim06tVX6vTa4QcFrf5leMkIYc64rfp7
XDkhEaoyXn3uI3gEEmge+T0l6Y22EIsnCqIhiBLiUfCd/aZv4pDGXl62U6pqSNR6Ph5P+Dx2GfyW
WQN/D9G4TilE7Tlf+YthAgSG6+RlhvB5atEy/BADXyDPd7S0BidozQB3/BDGTZVhbwDQssJ2xGpv
Mv8g1+w2NjxoVM71ga5ahB4wVG8+3qn8tEpKJR9jY0rJLAnsFBcVqToJJpI039KGZwCK804WHu8L
IxFNJvTd90TKSTukKBOmQQauPW5whUNemoZPpxrIH1ZU9UWIKFV08Xb9Vv0GjHbfF4MrtJ0HNBlg
IXscZxxSzl42Fd+1yuWABcRhQT6wsMEVvsitLdvTAMqvMWxGysbHYXqx3Q1WTmEbey3BQSo/jfrD
YGlIHFqzc7BJCoqr1Xo2jJFFzRJvjTiuvn6k+fPxUw0aKOh/o2xlxzLQGVkScUAkj0SBI8u2RWhB
IhMXYktS7MWI/BqncNlGnAErSo4hYBEsheWuZBQC509RNELkypTi+8JNBG233gH06BarpkIe7OgO
eSWGgdHkfQbTsSYTzEbW4zxi6OxazHHcXC9gFQB/vcu7uFnWFG88N+uJeNrXZRpLrBycaTUtuoUG
15AmtyQvVzG8+FdyLC8ZpLrQ2VyrIhMo7DdY8wDVeSqYSTUOKfBAomfuI6aaoF8Yj389ATVx4/BA
UacSP/Z8KgkFFpL1lzwO439yuIewWmHOmiH13d+TKYxSCrz6jqtxaN02NG1yr1rdLLxxNk1iD4a2
SsBY1/csPcNuFjPKqtzaWvU+wFb1oCD1BXyTyU+DC5zT/1JF7NijcmhClPUEQyUNoCTksTqMRlsj
454GBcMdUrWRhvvnS12rETHw5HL/CfjrRa97r5MBgnREK5QwLTfnLxeE0JoODmeHMQtsLBjQvGg0
WwW7sCUyR5uynFjprFTo+8clnvU0geA80NgwTSk4szn3R+NA1B6hNq6Y0PeOcLncHKd5VxLwYdJ7
uVBn+BIECChmhpK/fOdqCNGj3PBi+e8NRlcryDoOinhBSFxnssy3ro/znzGLx33s9dDBm8Bt9H87
9j4WL+d5Pn0J0Xzx7SnNSQN+CjYYqEp0o4rfs+BKXvjWhsUSq96V7DL91A5a6L27V/61uXKjOoKF
xkF/L7iEkpNgIUdfMkDPVek3Nosb3C2s7wk6p4NMqA1Qsssv06lEazhSI5JqeC4jbJjAEuJD+X1F
FmKWfpjuI310ZZGmMS8qFjsjEdwpUhKQYeIbQUqUJbm3M1DfA4GNQBPQQ2CAs5WQ5ie5MIDjEUUA
BDjWAUbEqRPAfPXnyB+ASAxEXFZVscvRx3w5LLIlNCS2sPpXEYdo+I4Lrrjy5qz8jIZRUiyIqTSm
3IfmqjXc3KS8mbHZlF9fF2jz2n9KH83SSsnisrqXNauAnNsnd7AUNHdaRV9eWPjd/Ib69tK0AJdE
Csqz46t4jLc16+zoW/bdwSW3wQ6gCCmJDpAs2tmt47h1B1A8dym5E5Sxjn9eH3Ooa/pDDlkJ2Z7g
V/sCYH3P87yREYP3RYRCW+Lx5hQm888aHwZYbf3UKYCsVnHAmaRSJ3shvVR7H01Z6dxnbb0AGP5g
LJgQFdYfDOtkR0MYvhKWh7jwAXjATz7BT44M+4WHm3L0rHOSZPbLqsYA3YOVm/Jp/FYsQndERuDz
N843TnHo2ys3n12ihYSKo9gHN1N9to76cqDlbhCpR5HOEQhxR3lp7xkyp3IZoNY0p/5ZEKLdObvR
995GBL9i78oRYP5bMn7wvTPkWErNmhh9cxJB6VLk0313Ks7Cd26YRwTNjW2RMxAb+Yn7Aozdoh73
ukMAOyTaPV5faVxaUzd/7bc192IcR9gWxztINi9ieJFT6QuQOzcK2cqjQ6aYTpZ4/yTjlpfp92Ok
Nz6weNMD14GAQDBRedVdZ51awxKPzIT+IM/DJE/2Ku4RcxZbjKfVT4rwEsQG1N1XV9ISd8Zrv61J
nDZS8wWg9FHkeCZWj5eKgqOEwHJQO2XpGd29Rf2oCNnS3wKdLgibX9KGcFKYy6ikLbFMvoezFdgn
DUT7vHS+EZXtOA9qiZmQ3mR5efciaP+hAM69UOoBbeX0DOj7QZ4jjV3M0r8/4bGLsqeVzPuhu2W4
RJJowaVd2/6mVZFnueEfxnwJx3WhuDGRMsAJmjhzE8TaGJE3Wf/gSeyXpXbmlVOzqYeVl6xZsI6x
s9EhWSwuJnp11dnLXWiumj5lHnZ6T+5QYeL0MwTB2Mrs4eEk5umkuvGBWr4UOh44tQs2zMRHHb9U
D6vA1X79nsrrhPxFyESXwu/armwGdvnZtcKRdocwrYAizEBc2YpAK0l7LUZBkFQLaglYL9aBDdwN
9Vwfdqg0GS6LU7h5Ena/wxVxGVirOYPMhx0mLkGYI/6pn3jMLIWXfzGIlShlw9GJVMHxl7A6OAPF
XuY3SfLdeSrEOcGe7fA3xnbe6b784mh6f0OzSfWMKsMHnWbij2srpSL1lfz6lQ9YoPPvU/MInQp6
OMmcDgG+TLEsqQIi2LHQjawHlVoFcB8WVKPKKE+PImMdxSIxHsati70FBh4DaoPHLPWTcGya/a7p
bY0oJ01A50e89sBjH1F/YUdViBYwuwxyrG589OKagPSX9KbJ7W4XEkAtO56Vq8YgsVS4nLugbgHN
joIYYOiwcbBVzdo6ZUfpPFafctIyh7PLhdckXogbWcJxEl4ImZKME2IhxFcT6ZmeMr642nvMpa6T
QjnVrakjvUDSNoPhup/EEDOGO+w4YbVFX9hDsgYboIv2U2WV4/afa11IKrQEEIIMJgSofC9LMTzk
+MkMzeMr5lo4DZKmYWoa1iKQsaWoJWqk4siEWM8o+GqapLZD+sQH5HpfaAK+SdNEc/3WOmc6S4sH
SCCoEm5PNs6j8JEyPSLe48fSePBS/yK/+d17GhUhk5ZSxpYbzCWz1AuQggJiTfru6ioA+w/jJTT6
mZtvFf0XB29vcNUHViZjAHMt8s+zdejo+mKiUWruROXOOZK8tMb7rtsEAW0nPEPTWdSvKa/mOyW/
htzMeQH9gnJn712cEBLfmte7dX2I5TbFd/niwfSSqDmSDjL43fhLOKo8Yxg8HDiXiLWjSuqMfmnv
A4rOJ1MWNRgzwBa+tvjOQRwBDbJwyFDcFCG8iO/5BHu9zYYMgiQLQaGKd7+2z8reqXg88sLgTxyl
X8O6NywunsJA1w9uefg4a0i9z8TAmFz7QOYuN2fZRhnIcEAv2ZjgL3CgNewrx/e/RrPdbwLOC0Lp
LB/vKNY+bN6c10+WI1xGcWeV6AaSNBjP6AkGpUa29bLxHEmufhe08VOZqWuZjy3qzld6Lzi8O+8l
aVKMSHBVnrNRtD6tFyTylBF75Al8lApb8LBLEPGIL2bfL8cu6YqLFZDcIHkFOJwMS3qYMcBq6EEb
1uzmkoCmD304/L888Q6wEeI4bI9S5iCvbcytPz0XP/h6DBt/13G10hK+Osy5b0AT6QUxp2OzkAju
yTyvF1qq7g2KI4yMKK/ePVJj44QzRWP7QlR3bSl2eXzzzKCIroJ9z10nGWaYBAwcmQkWKVW4/9YE
clyiRAp4N7w5nbVmnY15l2tGkGB86IvS6kZsQanBRhN7vLqul7Im+OTGfXNTmOvEZAgbIqCTa5Ry
6bx0q/7vf817dRbsfNGX1yrqbRYVYSV0oNCEMw/kTkVZy8Y7sU7jGGOJrSmoXIJw/g+81xjoMSIq
CqyiunKoRvDGpi+dPZq2o4IzYUjbVuzr1bLQzjDjF1XqrAsE6wjC9cnxw0lLIk8jk5FaE1rvaiDd
H/Wan5m57ypEfxC9RKTsFp2rfAF8EWpAJHSA/Z3h/O7ZMChLNWKjRR9vAdx8HqcVybvNzaT3Ov53
565LCmZdLY6P7WfYVD4TkBOIcqXGUJ4tHPlP03hxwk8ieu0m+Pm3lNhVEofjy3qRyzOjX8ULk7Xd
o5xfcM8DxjwV8xd17w8iSHCM6ZQrcfM8bB4mf8auSZ4f+TArT3+lx/0aEMvFGCChl6/v35kmISJ7
iPDZtl+Rc7pGFQJ8dIKkpAA4Mcmq85dxc8S8wIr78GiWq8T42/YZ6ELjeubbqcx6qNIUefO1ykfc
Ekr798g3NE/TApqoJmfIExHZEmjA1Xv9FfFhG87TFOGawZ+VdtHcagfrjYOx1/jw1uv3ntLdyZvj
BxZTOJpBNqAB+/UwZhyLFxXbAWcu02z4xQ0NaoZJcu3t+pHPlMlSI96QpZW23eFttYge8sXemDUW
ZJELvh+LQ+rGktd7WxTC53l++fmdagaqnpFQ8PXM93z4eyTwuSexeDUlOMYIJG4yrDsJzRZFfSkM
RtTm5JRaTqqCFiJmDwVcLB8XZMDwpOS9qW1ApG0f6NIS0NIY+hG+5Ul/mus21OyIhH25u89w+w59
URXPGlbHyA9OOhxWD657CB1bPhoM70g8yJCeWtf2+6M/mEKK/w/yk2W2oLHSVfo/eULEDuEPwzJF
jIR6VGIrFCZW4KBCtGyxHeEoaLQxGuqSdlQZC1IwkClB83/JZMRvfq0XkDB7BEH9zYZJ4ZMpjCRl
OYb50N2fqQMP4dccQAH0v5koZznFkyKSaBacT7RcAmdlHlL9jrKdyelkS+Hsv6bhEXn3GDAqVdsx
RnPVWMb/eiQJPzrMj/HZILzCMFu0+FXwqXVQ9e1P5Q5uGxlLDFY0spyOkVHow/u1Z255zQ17M2Gk
2KUUfh+jkz2Z6FrSd9Cmm/lDwaNPSOsptH3BmMU8gjHWy0RNqpWU4JNl9w7nhouLwMroo8lDik87
660Oh7s+tsUkvFdRtw6pnupCwpW89GJvHSYmF+usPKDvtI44fBMzrLFUBJauGr7uSVb0ZBTw1Nw8
+JF9t1e9fkiYedL+tvzcnbmHYI2brr8w18DQUhP4UAgyx/ctsqGorgLmkXiG6AC6ZOut6kTgjjn4
5AYseg5B2MVVpYvbXhHcv+svO2yZ7Yjijg+xjQLZ4s21BV3toWjomBBSQISWduo8lSR49kE7jMqn
piZT2aJBg536JaEs1JQgQxgKxgQZ59U0xXCcyJmlMIlpXhLFSkPba1m8WTH2nFQb9z0guaYGwsvB
SVwBTQkABt32uxxPvxwpIbf59EeIf6r0I+Jp0P/s6eggLbB9z+ZLdRWml9FWnIRR6MPjBWs3nkGa
5oiRr9vCeW7HMB23t1rOXop+OVxdNy3U+BAWX8qQBYnRGTPPkuwHJdyIX2Jsa8reahjIcyHJB7Ix
AKUiJ5ArkslBLB/vzbsziRl9CsBFxj1IhNFzbNtNQlE9I98PtXOcNeshhlDbJqb66H16OidcDEi/
miS4MuJuBp0oX2Gmu2HhTYiejRhAk5afS36pzqdKQVrgAKg4PLQvvYKFY3qSUHJQ+bHM1yDjHlKx
JoHo9+06QmujEEpbSbgVvkxVMJVBcWjl2w2johQwfKAfsEFvK5p8VRshIFj6jpoKZFTlSlvysQS1
yVdcHDKX9Eo40eVL8Uc5viCFnsh6AtS8ckKVppqO+hTfP4LnBi3nDF5gNaKV9g9oiPWxb6ZyfcwN
mVCfon38vdqhRNsc+6vcpQfYVSHkgGj54E5TtsoNUzyAnagG6uS6uwjCZJMTYcK+KrB3hWOr0dGg
pTIdn2wM764xGkhuO0A8meC9MVaZD6qfASEFplVzdKFRXY2peszOtyOZ5BNc+NSueF+//iYPXv95
VwmRLdRcrcNHvn3z+6xzD4Kmh1Emh4jcQUCuC6gvtif+/iLBhndQOvk/n+ijsHk6reSD8MsaB74a
c00uRjW6Rh6sV/VkaXoMvPMeQYHkgy4obVBrzKSDIprenPQVqvq3B+kVeiC+cw7zA1dBUPGbH5mH
/6cnmIwU6wZMgWnoBxfjIUkClyr0PqBjB3iFGT/f/8GmTpSdpT6LPHGv+R/vT6sVy2Ryr9dqblia
XLeWhTfDvLZU4s7DKq0WSid6JZZ6rMZPdjsWc44kd0jfzXV4PuTcXfJ8kv8IrS8wCSw0j/P8ijGC
Qp9ptAmvjAU7suBhstHA2TD96BzFK95ACqie/WKrUA/MkoZ407CYKTfA2FiR5eitxvJWwlIpshRN
NxLbbvQ3JxNPfKifLMdAwsVeTndiEZ4ZGV9DrhsydDWIyVzddxCyP2XuOx4G1N6vJ8nCiknBZVbV
u+YQVj3rdbuLQ71sscUiQ+i3mJ1G36JKTVIiGQNO8aMmmNDqC/WUwoQ72yR9I0knUYNR9VhlaxIJ
5wKdGDtcB4kP7tzrMmAmtosvu4kIUTU09Q6+Ln1yYmHA+avt2AKR2Dhnkgn7Je6/h+SZQy7lK/vx
qjoUThWW9939ZY8RZbIWC3FIqa7/1hqb9tVSdT9AjAITGOELw958oIOuf2ng1Bg657uLPRf/O83b
CYTgj2MTfHW1rIrjHW2nl4TQ84x77d0SQObv/ZpxC/awQRRgcxv791HUmYV/9g3IvGD0enQDxGeO
WF8ilpHrmy0jDePCJyOrP/0Zf5e2NQ8TzLEF28eHgm+t1YY3vE1z1zNskT+0Fjsn2BtMyLk6pN94
y8bHZNN4p0JZhIZFowLTz0SDsd5AbATlmJxxR62TNNw9+6H0TQV9M20bvX7QnWfe34warNP47U9W
tJTB571/ZzX4MJ+/VrClyJyRwchQTx6ssJJDbXs8fRxOws9/eMC/RmZkfHRYp9KDt7o12m+kNPKn
oe364Jj2xjyIpDHnXMGCmcoO+zBQd34SrL66vDixFmCBLHAhZye1mL/0XwjEGVPZlMU+4Nx8AC9E
IafUAE+HGUInaEuh/bR37Q0Q0en0+2fEFyzLbGRFB3+UiaZ9szWG8oZysa/941Vi32GacdAhbPb3
2cbroLi6wRRhCSn1eI65aYJWckz2khYEm8WPRxH1wRAYfDxAhC46bM1G8B2cDmTMWm9rA1vC5GiF
xRGUmDkcbCm5vFuWtOZNGe7C7yagsHBE8EoU9CiVZL5xegwBvatbWS13ckRyW7cPUPPAwm7eFMh0
0KXCVwCLTFQfbqRdj+nRqcgAXtQK8VsOilk2nfAkXQsx7F8nHkT3vWQf0UUjNe2zOlZf19L8NXq1
NOO/L1dKR0CjCO8yEE+igMpvXkL5lQtJy/I8/Atu3v7E517tjm8QvVjYF2dZfWZCN+4lnTB66ZOK
22vwEOVT+HsqDHfJRxOb97kiKEuoPEFe7fIOFQqQlCbiKYEM2pfx7P8QkajRdzuaHcNP1WQCa6jE
+JRWZaTBwsbKqOKYsHST6GST4DfudJFgnjJL6MIl7QLsrfWgqGD5szinw86bHs1Nt5d6zWodUc2e
SIcXyLZD165kIo2l47NzAZqkr0Y+iez2+6oO1riT3Q5QD/vMxiuIlEhXXF0Ok99k4L9cNQ+emROP
pcxqU3fIKRfiVuW9ev+7XHLR3iZ+wufH+fKExrdAJPuO4f3FgvsEsbkzLro4TO1EKyh2aYMFGeDB
0D9XfiYlsIrCqKW319u4D2/XHmx/CpbJnsLDnu0ppS312xhOQV53zrt4ysJ9FTx0AFuP+hUV48cZ
ORZO8Fl4tbBLGEf5uKGRL3snufS1ohB9eyum7YxZS1cyT6BTeXBK4dAylBNoOpHMYeGvbLAxrWyi
RsWPtmnc556cflFUaqyJ4TN7UkD25FCqXmReY3/dLU91VXZvFfcTBzA+2lSZ48D+pS3orMHvk2zW
1oS06beB/z9Jdw5K40ZJBh3OTzCp81AipuLpMh8ejL+LsKfMLSxnXltLDd0iJJDWSa6/iBWp6DZN
/XeDy+nCTzKDmWv/4H+rMd4t5mhbDUZ4WNvQf0tTMuJ6otE8H8Zw5z2OB9aVpJiyJsN9ovIEBoX4
q5RLiJhVIZVNgL8QJE0Le19yiEog1iF0vcuZl2t+h1b26HHk+FUDTnhX+WQ/oXEAvYMfZamedbEz
OHWznNG9W7v/dGa6GJrpGsreStisanFNe/GdNZ7pxESXiEchGeQD4ku8zfF8PMMIpkVkkzlTZyJk
DwO//eyQyXRtOIBH7RksK/m/lfVnMnHT2H03/6pvV011PlAwEUqiSSo2ZX3kOLSqRZ1kdr16Tc+I
ypjBKwczRrrRCLqZNGXfZFP0O68sdqc2nSOLrRTaz6Me0wnY7RATBSTOe94tDJoAVXGGsQbdOTY/
zq8lJuM4aqbGl7va6i2w4Oosy1g3EgHYcTISRuSD0kM87zyKE59XYWJxJhXQVRJyps7Y6nhhA+UO
Iw53KrelTSxxvakX4Il2gkS2qN3+GgCswS4SclQ5GPi1TnzUNwKlYybWN7WpOtwJ4k17AVJB5aZe
ceOXVTAS29JOBKCImcIC5aXfTYhmmaEOk3Pj4i03zskWlJdqoBDYPqYniwhdRd0iNwonSU0uEeGD
If9tQqAflOasKRFPolcZ+8snND1sma/L//NzvUZ9kvQJiUS8IzUWuV8nLJODimz/u9uIFUmcP/UD
y9HV2SaYeBg2YQJErRFvIKzdVGa7muv7K4MwbbZ2n0wwO0zpI/YGfF1sMnssZBmkAZUBvFbURnBv
MKbO7KbqXFz7jV7Mzi7yV1T5UN0rqB1aYlf03AXG253MC9VPVDVcgxA3+mybM/bb+zfdoLKPJQMR
JWq8rKCbCShKW62ZXBckbfd9PXszwLrLtc+jyDL5zGhx1vtBrLXJotEyGhaDrOyrd+YoqVVhrIWp
QXub9aifcr4z9pS/IHWsPNVAJy1HKfH+zREUfmGJ/kJd9wqJVnxdVju9ikCFdPG96U8BgNLnhZZV
If0B/cWf4uDBeX7s7Oe+GUVDk7GgRvzDARAZqsybE30xjYqkFmmcL+OE/SoYZWHOK1rkTPUSfLA0
qcZFLVlP6aleBmrjiWcH2Zc5yRYsSJz2UgBTMr5AsdcKfEkooYVC2w9+Mz8Q/p5flCVy1Ye/lHHU
lqgp3hj+6e2ntRbuwY4ezTQR3B2Kca0ocJ0FMwM4elUxtN7ObrhUKD2k3aVdg2xNPL2zB3Q9j0vw
F1Ca96alEb5eI12+CQTBoPTNn8OU+fju5C99bb0ZU7lG9bhZtgNZhGs4cH5WG29GwnZXOY9yMxNN
j4rzv4Qyq1I68O6OS7amFDQBcg+RZlvNkEMZVxqY8Tj4glENcHxIxhQr+lTPxYXmn6lh0H5YPlQJ
TSkAnbAOacCUQF87RMOkJd+SpjxVo0F3ipKzP8+w5Bt14Wj+9mRixs5i4bma8T7SlUdCFpHQLv4d
WqtvnU94fzbvuAf/AVDAOzaM/36WccQZSzC1Qw2mwBdWrpuCAiXS+Jz52Rk1fKyxJ4kryAZpvJ8I
tAi9z2ArDv+AtveP+H1/bWbr1tKbOdZRjUQyRskoHhIsUwc6ZrTSzcTIRgZEZzaB86Oh6sb0zTYq
Wwxi8MyMdilN09SKQw4RuecmD7KMeEav/iMOBzsl6rrzRlLYIJZov8y9E4blmBrAWWc5mtEb86GA
e1EdKFvYBxlFILVzSLFqFkablo3mtyZEZdUjTBUArWIZN0wnLLW+llqk4psBi3B0pf4TjZPpKV5p
s0gDciC9jw0q31D/qgvrBB6j7rjc2qwkhoX258vlL1jMSerXCqP4vSHwjWNv0r12YYG+GGsV1dWM
1fyZFuMI2mPWOc3m0fxtTiiJdvrKFj52XxhJosEUtGtoNtrGWu7DLScTP7P8kWCq2UwHd2SEB1ba
paIEcUX2+nJy+qPILXzEBwqfYS6zOw8H5AEU0JNvgHPNjBSzWT3cK7vAmeql0oG7dKaESCubW7OF
bu/BgcAPobxrSwL5oy8DCXjbQE7jndDuscWI6Q3lLs+BCHb15L/kkjETVPIsg/NP6v1uOJdnhXOR
rFjnT5UtVo3Id3ePmdhxViSPXfnIpZpF2O/ZPIkIWyOjZ/tWLCpD0NBaDZ/5LAnJIcwsqfsSp5RY
tXfq+u4kL9BdQ8qU8WJFrnwVmm80lyskJlvQPr+hnT1UKcVsJJAreIwiYQXwFFL2L3djliy3UwVJ
leNz1L2A1Bmi08aw69kql5rDpfpRUnkifMYFkN3YznsEpRsAwS8jeGWLUcUpm3cTQfLN550evn6I
7kExCDPlbodCPh9+WZEv+zBFF1JZHK0XYHOsmcj52yi8gr+qNlF1YoC413AgewTRSBWaV3Rqk/kU
DzI+thYkJBZNo/P5zNS41xqjowEXLjFubJJLGD5PXNb2Gi2JsH9pqVRmYOcmIDabGb9nmN97mt0f
3cO9yRm6tmsN2a5h34EH4luaCKNkoL993mAA2nfKdXlU2L8BQCBna5WFZl2CsWdci3SP9idnLzdM
FdXFYwKhK5/wgJX2VdSBs5QfK3t9fQLjo88TWcd2/L/m2c4MYIxd4vSHKX2Y+Pl3Ewr0X7CT+nUK
ObSHuRGllgqM4Mjm8dEJx86IuREsBWVcXdOZdXfxgJqKpG89M0fPZfRAfXtd4c+pSym6IbBom/6C
1mLuSlhfD3dEige/c6Latg1t53iZIsMRzQ26CvDnlY4yCdEjzZAJq5Jf+dyfFzGU4MJ2bfAdKiEc
pf+he0HGjVnL0gxyvPpv16+tc97ocTbo3WeaUNyoj2AOJIIQ+kIyKsh3J702ajLaJ9dnv6ba+PaN
w2rsaIl5LtUZ3K4SOUXcB2h45ulv3WCZrGMEADVEIMhX6ZeJU0fq6u90eBiBruz7rfVT1/VghHF1
S4xDb47fM8V4lB5TpCGE9uOdkXCmmr6vgS2pllZE/HMCQBjqD1H9IvSTUUaDk82i7qHJmKPxBniK
nEzqsAqUrA73aNNGa0WMDMvPMLLFfjN4UNVzeeuaXjrCVwgl/0T7f/CTa05OB5whhgCEfca3rcLN
bp0vwXGHCW1ThJMz5kq7GIKexqVrGb6pkONhtE9MB5WmT5xFX5Nst2JPMeDe/L6O/4hREOskrxIu
0FLscLS1pMCPscYUKAFA0tJoD9MvMS1tjbxtO4B9qqV1nEaChYHXCNqwSjZJisQFIW9hF2Q6UCTC
V13EumyyK0oc0DAxm0UywjRt156aZ4hzrw5L4UionNOuUytp9jdEmpb7yVUwCruaeZTXMNYhjv++
7IzRZ0CX1UwUJxoPqDwFl9+tAzNwII8AmvKdY3GETGEitRj9r5bsSZt6uA/g4mz3ELIJNN110hbp
I8z2EVTp+P3FmoV0DRK9S3UK5Y2mlnRKasWZdjxLRSP2voWdnkMBBZgO8iucW/hZERl3Ht+AHj1e
X/O9q3aefs0RtSWeINryVQHqI67PchnJGt6Vw7+rNfgHoLQ8T2EyZQOS5aDsJCECUlIJq10yydxC
L8nrB7s5lssx/Gz8tZmFHTiDKkz6UA+X7ZuzW02kjCL64LKp0t48UhmDmawrUL3ycQVID4yi8nu1
LmrNsmpMWP6XYz9qb18qKcas38/CMEP/J++W8LixDQcYoBe87GOaBd78xrMhU4guzeXOlI/V+ahc
uvtOpB2abWzXrIdttk4UclNIL1Ptb777jGygnEjArKBhFdaVsQ6gzRrBMvZlc1yTJ7t7bR3pN17t
/80cXklhL4+oxi8kJznLh6+EZEZkgqiJYulO6z6N+eMb6Lh8BRAIomHN/6CpHs3fIX5yj7oe8W3n
ADmzlsHXwPNilfrg0Cb12hWHOq8KNBJNCCZ23uRva/Cd0TpJecDxwq+11KdFtrmh75G/KC0sq4Ym
1fqw/c6BNTPhvLt5g9KO0vWhE4XQKxpZl35h3OMmnLeV/Q9X6X4l+BzBBE7K7r8/Oz/z7vfTrEmG
XYmf/U0iFXknPjSIymbLIBg9QQvgOr2uDI/7ujVliCRwWiURM7mSZtO/4Ebs/uaD8pukszknn9U+
c+EiAuu4yKlDfYXwZAZFTzT8jEFpHzmogm3zunnZ9M20BeUh38ruiKIE8xO6RIwaXrVV3i0jmRNE
7SxSDhty80Ia/zLuVl4hdAYK9fJcpbeOeW74ql+tNHrhykSoUhmfl2puaWjTTLWDGTRjWDCRNz1+
EU9qhPg0OxF2eQZff7dDw1XjulAlAaegqf/g3CCxHzHoUUWC81i4wmX/dIz6CqrtfXA+rrnhhkop
YilKcbBcDzIoIpEWXvwoZwj7cyLQxeusRLxUO8A3QFAR7ZsQBsmYsQJ87iq0NI/J3Yic9ZeVXXdx
zfa1KuUF+5oRcUQVsVJD/hpbGoIr5hsObh4bZ4qpj4T7opvMD3ItHTtAeU1W8nA618BcmNYCfwgP
bF9GDFa1r509HxSsYZi7ThgxZqCtf7qlS3WWpeZC+3w0unlod07VJABj+aspDLLaHQDrdZ7sKfMY
XddgOdL3us72hHv1JCxveZznorCkeEAUCmS8IAvZhimvuLdzvLA2WIyncEYzkKkbf4wnnnxEWsBI
vk0gnAyAt2jSDXuHA/XtnLzbHwsm88Qs/9l2XGs00hnSp09F2HVI968YvexS8TpOwmcGDNt1vcCn
aqUwujO++HBvYWTraRP3VaEATS6rJcn3N5+3qGiG3BwTMwAqoz2AU2DPep+0uQXYGyrGFCyNp/u3
O7JxUqTEJ7NZkvWguDIDS76JSm/wWWNCoCjllDErR8hXNUeAEF7yvaoMDR5rXogPeNjv/X+joYhV
8TRp7tKDa+Ogu+R4UT5VlPIJdbJtU9cb6VOQ/fURE3jRJNtGr7+61wcclpCF0VeYaA+GBIsz3LVz
KLlAjjpYZS6PXldwDN6ksSjJVbjNCwGuVZu1j91AF3KxUTqhkk5xW3HOYa0QECVjlBGlCwk4J7Hz
z7e5sqaIMBxFkTuRcLJMuAZGGi/ApFbS47UPDvVvKuF50FSAfkfPTyK0Ih2ndYc3OdI6av41WVA4
RG/3vBHZ2InkN7IKZ5Uf9J9M6OyA0nwMiBUL/2EjFE8gtS+j4hiRpsvqsUbXw83nzw7rTbvLndB7
1LZyu88eZq52NYBW6wlM+u9RjoUQMrpy0v/KT5MHyVVF9nWjg1AcAgMEm6B1IFxV/9os4vNImJPg
n6vKgGKOl9K6/n7f6dDd9J00QP+RqdjsvGoDD9brEigQu5jvxqKPrJUEuTZUPQZvBJxKtMTt6RxF
sIjLfoavF+8kX13br51srh3ywSsbtQwvFFmXuL9OLE8pUTuy81sBrRNlm80Ev0WQEh3ViAvaQgkS
MK4WiW67awA3UeGnFK4OYQWc64xT792xos/CI+YrzEGgZQ+NZZVw2ihLxcQe0J8aNWNKby1xeK4J
9f+2UDVcu43E7nyGZ3mDSp/vyVnLNDVZDhk2n3zcR+PdrwkRQ27fdtmbFFmVqT6bXXFJanEYxdX2
6eBWRvD2Gu3kpTE/Oy3VBUKEtiBTs6WhhpmWI5gE98NZco2LU6fdgBxK0sp7BuiKO3hG9dE2YT3k
lgDPCvAu1eHFTm12BSlYMvpOXvMl0Z1cj2Tqiu6FoJnhXiaLky8F0NT5S/fkSK12hID3sMBLd796
5/Bz21cUXVf6LjFYfB3kYEo3Hbb4podjP8nFaUrNgtuAXltyvHZMLhlhPTJk9rCAcpiVrqGaUWxF
mnmORgbeZnzBJgt38tRr+gtOrUBANBNBm5qDVZnhxTWgTWwmW4rPtwzw075enrTQW87jCtq8Dbc/
HxYjZ8Ei9b72CWVB0Zmtpdo5CSDEyfCUOc8tY+609f/Ffy2CP0PC9fdowDKymLH6uUDBA53gQQ4Z
03dKcKjwWk9+WZ4JSLU/T6jlD8R6681ZGBkYjs8yQBgqmRDnyHZWRPGD6xu1NFZc1dP/CR4mi9en
9C4mRRr0ES44ExOxBDk1JyUM7mp1OqP2Xx5P9mdCTmUPg38DW0daO3ghh2okG+sNH8SA9hGu9O26
rEpqdUuHrlcJY24P/NYbcIQ5FkDPHiTnRftEehG81FfgSKINYQJcUu9YhINWHqf+4JwDuPPWqRFB
oP3VQkmCgD8YNbBvOoGLgDZZPMqokxb+4/MXW3F0dJS4ZWI7Zlc0dHLVSDcukF4rUmlsQeWxGm8I
dyPOMjv71AtlqORcwm1FXZ0yI1yic4kAxzrIUERlkzVvQF+IRe3j7s/t826yePlstm6r8sEiomVS
pW/0Gs4GCf8dPjUJDV0tlMUjDphUjpyVGzV9D5usOQGre3STxdvO+1rblvajDzXTolJwWwqiGgry
6OgleIhjgOlvb5aU7+Ps+DJIYtgmuUWfQD+QvJ8BbtGlDXJOIbPRB4esIfwCiK33hqxPBOVTvus6
AoyLfDq5D2jc4RpyQnhSV2UGJkLm2QH7T4+Z023GKmwoz2BPQl+Egr7Dv6xuSxHJ+0WBJ3Eri5Eu
Ua+Y3tk4rZv5hT7Wx3jptSnHSn2Sgvvoloxk6k5RND01JmqMEjawiPDOURa0Pd74HmCadla1F2JI
oVEWwWwAgkMch8VryTc2m/0hLOnwSwSp3GA91E2piJS/OtqCWfROhBJvq6EkgEJB95/jDjDoktNE
oSXuUwEbyhMRZdAfd6bUnJU8vNCm2XlHhR9W+RxgXICh6FBXDPWijln2Dkn2aKq2g7dmW7ki6G/I
N0Rz5LQAa/ArRXNqb3x8d5hPT8DKvgz74qs69FY0en4Ywj0K3IhEFZgAPoFVHAtiz4HWOrf6JmL/
ntpp7IpnQJ//+Y14e4O0q57Uk73t7L1bkItFhK8m3J05gf6gaiiJ/e/F0UgKPfsoREhRDI4npotA
n2yU4OqVkivlsErJokhilGPd2jWYyHexsZ61/gbFLROsxmk/io6zFVvaLuFJnoLScFXrmidSYFz/
nuWG5viATb+hZ8I7P69tDuZoVO6W7GI9aDdlzobDZylHiR+NwVCPbwJ1QR9uK9JcOGJZ98bQrf8D
UGdm3TxmFliTPn8wt6cCb71JcvRNPaittriI09AJCkTKlowtoSql3atWfkBMN1ghNx+6MCti6mge
y+J8pUeHa0wO/JvqeHbvVbJi2U3u5L3UdqKpAhJy8vBLSidWQTAMpQxEofeN1aiRa8ZsfuYLti4V
4OvcpSXBhvosY/olNo7PUcM5UVlYi7cRJWSqSSMAoWqNuoWj1gtT1rPkBDvHFdU6XZG6RpYfQk/7
hmWKFfoMBNwW4ROBttW45edJ2QK97Xgz5gd4KgGI/Mavd4QwtEoE+X9arwtuHx6sS0TzzMZylSJP
HJoMxBbO1minbSskImTN9riQlAJujXfyAQ1dBpvz4v5ftzAxyHjRBTUkZjzkaRiL7okltJeqEwPr
vFl8EcYcQIcm6bZFxJCJYWfvF/M+nOw7Jlzu9+Q5d8h3lF0OHqX02G8EmWKFSkVcP+Ff3xVxJ0DT
Rd4iqa79nVjJXHIBtX0v7eI8tbnKVIaMtdrqXhR7PMyKUGkpwXo1bGYMLzrwSD3KtBAy7ekWK/OJ
8NM0+ai/22wmpOv9GrXgpmt3Jvvt3+clpvZC1wOuFXVgNFg9IHtyJk/yTMtzekWDj3oTwNqYtBE9
d/xQXub7ZQ875o0MMAorF1BrdLJcmLbIG2QZj1b37rtiB4Y0u5uGN8/ELqr7uwRlYZTOcfk5B5Fr
nQrNHT+v8ntcAIyEEIWTIjD+OnITvgzNdXVCK249VQTZrM5G8DhYmGl7RMXjShXDBPjh/xp5uWxQ
mAUneX7rJvBfk1E62Q68nh2haHe4Zh2qprdLAmmyztGFk/byuNtO7YYIw/yezDlf1mdj3pwHxPiA
ujpDFOtzoAiT2JD6KCjTWPISnIMGQxFmPj98hOWgNHyiml9Bev811LtO9oxJlxLnPlTS+jVqmqYn
nAWfz+dQSGxtYPN6LzUCC2vhb53hSCRgkF/7usRvAUVa5QuPQHuI5P3Uw1Bt80QojmZHF9qeiGkR
mMcY7ii3FA20wgRDtH0+eOTtDvzGBYuqKsbmFOFu5ca/z892o5Px3W1L+xA8MsB4cKom+A6B/ISw
cs7lhsXMic7vwx9YFjIlVmsnujkk5pHhQQx6ie2X6AGP1VA3nKDpUnuZlYWBrxVrOpI78wg7AXe4
a648oonK3bL9qH6hdnejrGIzZ2+yPS266gXaMO7iOwx3Bp/TVEVw1Y+2IsSYnfTfPO0Jbx5oqmWS
0/Vac2EYVX1mQHzLEyOIe9cNN0TgITMB6SdFDbmFGPogaa6conLYOZfupFdlhTm/P3kgI0IAdPBY
0G6j6fkVLS4e5jIKSy7pzh6ZWGa1CKntDY7DBBeiU0AVCIj+YXZyMHWVfQ15+0dfdYuCcPgOCU2G
nLD57hSwEd+ZfdDoZekwdGL7Yy5ZVBecpk3278zHRV+EjgQN4b5IJvZFnv3yLivL6paRKFjZX0H1
jbVFiHcyZkKcYt+PFcmyVDMy0/f0B9khrU1EXxv4BxZVvqhy6P1q5kE+I7EPX4ac5Hen/+WpCDwB
DplGPQrQ9syLuSbOI5gE0MVRiBt00CPbtCLstfNmUB4V2JFyT33Hu40NSfcTqQI99svKbjt4oqJP
yNae3MCwEh5cvCEOfML0kTfRKXKrEfkG3W+BUL5WWj93aVrQQJhP0AtGQLUqiMLfXdivLwP0bQMu
1xW3IzV9ySCsKhwixik3y72imKx0CLUpsKZ6tmY+UvsrnU8zMFQ6Bi2tUJhlEKudX1v4v+ML7hfy
daSp2yzw16wT7t/R86NDIfg0OIrkUhubv+ugCYl9eR228zAlJ7t1Qogdi/T8zUnAK+n+hTUvIl7V
ZR8go5qLE6sRnwJF+TQbjCT+Hy+Kb+LiJPiEtS0+LI1LLDKg2ktXcctfLIKeYZPQtnyPJNW/vA32
jIMe9dRFPDNTJf4hkFBfQY+1f1OQqqc5qKPPjaFELBIycvnOTbt8e4kTPPaxd/Yz8SK09L+XN+85
LfG7OQp/apngzPdXF/1E5JvtLdfz/ZRLKoOmPcuEU03c0WnsZG2ZSIe8ViIDDRH8wdaNfXHB/0nK
S7u17OhyCKN6WlkTzfK4KkAglrAYDIiKsxrOXDInQH9rnvTxEyRXPPPKbFhev7j+ZSuf6bgHEEKP
0PZLUzwRSPQh405DDh+T6Gj1OC/JD+6mF+h3PYc64R9tnHxVo15wMgaqkG/h7NPeRZmIjJummYT0
dlSmT1poyc0QmKYePiml7KPntOrybbVKNXBu8W7fYWnBFpDNUVDRj86vHF8I5G6oIPa6sPdf+Ap2
06I735gal0otTxEjQHrlSp+8hTsChTsCD7jKBIHggRw7zUr7p0gT8mtfmdwuFOjNesqx8Iqm/7y1
CKdCuAI+k+m8mymMG+OGr8sN7Z/jckCdLr2g93+enx0eOjI3xTJnqD/V7XPVO6ctcQwLruWz9S3g
w/12YQ13n+9II8IJ/zF0XDPnA9wNSKGA25mrg8nPgDxOv+gJePNOKy6NPq3CDxZ04Ou+1/ntapFB
E48Y+dW0ialOMY0hHI3tM1NaqGI4lGMwf2/fMM3vg1vt8u7L0UJi22c6qfZouyJSA16G50JbkQ40
j9gkxDc6KkBcNDJ7dflmDuLyjcO5cwf7dl5TagHeRZVRDcLQjvHInxXAqWZPNJt/qvP7cZeQUm23
xVI2JumoOITvZXraBNSvX/de7dHbIYigqwondofLJBCcJBojPVMQJ59Pm6xMBTgWZnpT/7lDR8Ab
GmBrpQy01Vudz146IGDobRjMp0zujcRIbDBcx68mAiBw2ivxdR2IX51Gk6V7WgCixOWtS6TaR4lr
Nt3GyOwlCzAj6jE4NlRDUGWPZfItZh1DX/mD7IumvTTMHEF9+2/ZvpeeCkkFRvSj4MuWOaapHNMx
NUBen8aK/a03ldIWRieVuT2EVAPAgvhZJz96ht9UOc6E6QjHIlHiyawY0iNzfiJnGyg0jMj6uG6k
EBo5y4kRE8L+/G//JCfC30DMd2DnIhqPwPIlsdDR2+j5wmTWSKk2NO7LqS6zsX3XFmir8E3p3y75
hbbZnRLbP7G2KbTVi9tcklFy66h+VmrGjcqve3vGEzQV6efIh7DtuqoktXm0uDxjwfVEQUMMPf+q
57oUco3LFUMdvJiDisW+bBepSj8jtTWE6E5ITMrZzl1sQniAg7/xnoObmyimqHEDvHF34TJ6eVku
57FxByoJU1OFqvuuNi43OTwji/yk8B10EE552IzaeZ0rgSfhpVgKXBBVmTLAiTTzFUbmaqMlR6FK
MRpfpoe4SVlMsrE7RqYZTsbI2icknloRmaLOz53h3BHTh6q0hk5TPpULWG2TcXUfUGSp6SAA0ONU
pulMI1Jgs6I83lAFlA4V9k+DLc2tJJccAFZ9DL2bGLrcgb7TsUfOTjthVoXakLTI5nM1jlaDXk5M
SNFUQSAz8Scx1TZNbw4WPjqYf1qcmvsKfdbxE8YIsRKLJrt8jr1Mpxco+FTykAJ/2ZFHVmVTFrCF
DoIPYhFkj18UzTcLNYeNOeJwHn3JZ3SAbwbe9SKgZ4XvYED3AlSWGkDxAW9eksrbPXVFfjdHP88n
zQAohQ4X8bAtmCFx4EAcMSYgb1x2AzED6ftftZX5SKJd4aDuUmr2arJcOX5ouOmbvDzcbqldbtDp
o7oFJghqOPLPTna2l7zll3tG+Ic8GQpmrb6xBREVolGgcBeXn/ZM4ibSvB9IWI7iXcp5vZ/ut8FY
Jo7DlBThDxk3XV+XZJcDuUSLuloSptEVOMiBgphhL0ASz94VP8kl8JUhnCCz2r7Jha2w6uit5r3a
veU5QVAZfloFhKeBtbiy/QqqH22swyUkwqWV6F7AopOj/cczboNbaO4MLxwZs436plMYpZ5KTLDT
Vx93V7idwo8pJTaxp702w/mN+SbKQLivvwMXcERLLAk+XTeJ9ayyU7COMPDQ4lfrIBTj6LJhUI8v
i4d5AT0Nk4lj7MEr/0aXF2LLNPGj8s5DwauBthd9KmWQdLb1JLfHv1p+9dYOnw1mWrdhTXT4ruRB
xfUTbrLXjiJ6vjzaDSq6i9+a1zKBCi7YO0i2CUFFfsg3QoS4ydP3K/OzpjmEDIzBb8mHs793SmfQ
W/aDIZenj04AMM7oo7JfqDTKHc/KO5ltN1fuiQzxV/js/vbjBv50Pv9pI6zhQF2kSRjY0cgTpdfE
U2FUbF30PAUBaw0KsmUayRuFOxplZ85vWksNA7zTe7tcG9kxFVCaCl04rvZNkQXnmndLI3Mxo/YW
u2qLyBtOseSKP5C2vnS5PGr3pzDNawBWRLr6Unirh2nYmccWrlK/B99fkLc0PBHqcmKnjbIxwP2W
rb34qkWas2pAuQPOiapEiXm4B61SGMQiIQc9PC9dzTXtn17Fe8wv35tx/x8QTaz61CfBabHeVKi7
VijS/6xT2uTq/Z/RzhK398icbIevgtjoNqUif5pNvgFVJyOd/ooP4HNszimqAq2zhyVE2NjtjFpN
awsWNNZAueWjWqfo4jYP/hdlxcjxC0fSmZAFnz/D6gLPbzGHG0Wusgfa1TQSoGP4U7JgZ/1l8DMj
coBC61uDaXf5Rl36fjg34veLw/wC7kyyHpcwZW438pNgtjnEY7w8IzWz+K5pxQOoj5rlNENMezY4
qvxa+dByEbCvLf8D4FwnOnhyUWYQTKRwcW7UdB3hCChWBn1WgedY/rAp2pIwbUoOq6DonM70w9r3
hXpgMDlTPsWWeG6c2ALKhMEOqwGI/vsOdbt0kEgll8tyXhwaKPHqUOOvEpDvZqCTh1ANUPwwWNix
l43IggZsGXUzaFKmMSjxVpcISiwyZwpjoeFCaeefcfhTmbSk/E1wrbB1v6egMOOx6Z1mRWTJGR4n
VwkGU4Fldfb7/152n5IoKobZvJXPWPcydECBLX25H+qD80111dlZMxuRykewVOqWqfVK3a49Cij3
hGHd97Rrx++u+HXGCDgR2kUxuNM72fPDoSKacIBbjYWXGR12Lgm9lSQQuEIJzqlpqh6npSq3bQv8
L3TaBXgc/D4VHHsFB0YAwbFNAUV/vLN7N8R5jOnMNgeyOYSY5OEdUjyUDAa0W+QTsiuUmCNYrFt9
yM1GNdkMMljiXDHVuWCaDwHXnXGOoQk7L6mPyaElnOFObkkgO6zb61NFf/RFan3dZtf5KmHphMps
iTHudf0gEgLlP20zPxWR4RdscW0W4qYYYkhmDHUlI3PBe3MVuEdmU4bSdOmJwOqFDdhO/NJz1Kdt
BgDQ8H5GG1J6IyeVj8MW6U1r5KRi76Kj8J6P7gDXWkU1BMBSTI8MktHV6kT+/Q7Q0/l54kUvG9+0
63g+spJL17sJRC0o036qQ08WNJ3Hz3j9dK95bKghEwH86HSW0Lxjx2CQGMwNOS928G6jDChEByS0
y5n60iUm4X5UY4AO6LJJkM6akqAikoSTynqiZ1nk3teMlEC7eYH3O1pwp27+F4t9skbF0q1QqQRV
oEXoDaYSVkinE+uB5VP4DaeI7OFLxHLevofwuzHtap3zk34PwpDIhYRwSOcMjPkOTvX4iwGKb+Js
FhpyE2C0jGTPDMV/trAXPHdYcqSslffR4Gc9Pd1ynirbjCYlzKpKQnTGiyH25NCJNra/kri556IL
tVkl3ZsGLbqiRRqhEbbdyekY8ATXHIpoAPDQru/yknO/v1zxEDu7yW6IItBA7NQoN/8eSf6FDzhd
hvWyyLueFpQc3nYUB5O6sljC3RDaQVb69syjGZ04ffFs417GmjP/o/3D6/hR/Rbpx3+sGBSh/4Nv
xzCvBlMb98heHqyOnck1ntnuaoof4aZATuapG1mvFqYhFfBtH0zrAUWLG8XzXgbeNxEBWgyWcsFd
JJS+TbhliKiwxT9KGsLx2GkV0YkiYfSOtvzUKtH/Tccb5VBusPhDZfLTxJBDxdAiT0SZbgByj0M9
5V13mll3QZEFjmlpuEWchCz1RqfAo02tQZN7HzczvBcBH4+QMpvGHga/sPtyXXTfRI/NuQsr7l3o
flcXSbaiD3lbNN5ao8aHCV0jzaylTFFyhPVYLOOm7cuIE/XkP1THQWpRfednQXlCH2EnYY1eMtX1
RISoEARQWS4oePCLswo2eI8uZNyo+3TD9p4a9enuQ3h+sBnU5pYOlgn7S3J3hoUgEtN4Ab9sI4tt
OEQmG64eakXPZmHLcFHxf+UoyncTmDrFD1lU9kzk1EcRGpWgLxR78z5HA8bens0ikxDQb9a2/9T1
ebSbPkONTP/hbaGXDq27uDZE9am68PZs+vJFcKOiMb2BODe+rL1aaYc/aIHgTluGVddaHdQlfnji
9V71ooZ/qrwEeScPSiZEKnYTprKcWIIf1zG8MI0CDiVgDCB7bzjdgVWxrZ4E5OrkjJQCfs0boU90
WxRK1oMY+ZGw5Oxwvdn3Ct74CEDY9BuqbBjEQTS6cD0tkuuPJ7AZEQEXQGLifrZmtA968fb/LDpo
T9WZ1QK4x2fwf9v/KZtOXD9HGRHak2Fvvj5ZHjyncNKGXEJ0VjWaHKg29DzMvfWikD5QiNH6uYA9
ETPqHR4uSaJv5wuycjchncda3l46/rJ/BZsPM2kmoY1hMCSFTqbvCGM8Don4Xcki9NK+GhxQlPcE
9PnXW1ETHZXWuK5pSH8m4qpXSTyeJGVs6YNIJ0EZNetg0viDoCNpVW/1jeOJ7D+/+9bcravKF0nE
H/fjKSbH6qEKZ9ELryU0oSGV10kLrlB3HTXbJfI53e/VWZinn7n9ncfnLbmIZu30pe5ST2aFTXI0
aboxSCw8PdXBR+YjjgIXR6jhHASmTNfKR3Gw33K+KshvWgpmCQpPuP9QdU9cHCkU9Sv5+g+xwMlQ
uuD+9XzZSIg0jxTg7PJmbUUcSA/R1FQ7rVPjYSaWQpe2EOv8PX1aKq9T0sdl8kIEnEN6B+qaZS6w
gmcIipmAKhBw01/bD8Oq01A/JjwZ1pVrLbMxtbVpe0+PbrZ4gnrle4jIMKYpsJulJZnhgPSaWrkb
S4ybFZqaSeMW18j/x5eXCxeNQvGH0G9D3qA6MsO8lF66bF/FX6MuiOUdvdGVlzErgWu0ZZM5OpVQ
cNnPUGZr+O7Cw3ZL06QnnnT3GIVzHwA7w1NB8TyfhVuOAms5FZWOS9DxkOqstsiLQ7H7nDrQkV0s
xn2jUhptcStILwhj9BxAzoMWwA6jT0X09GKuiGPUuk/q1W+qdHlas+66HTgj3FEYUlxrub0ypTqy
3IJjP2h8y7QTbawY6g5yGe1+6vN5TmkEP4afkOJNSJxeCEHie2oSAK7TaILUSBjSjViVtxmV8GGc
DG4aPWZHU0l4qTkHPTr8nIXJHUTqamtJ4In38sSCuuI/5QDNEzUWpMjdW7/v9PrfD6RIASoLZW2X
tJmnew8rhvcXDdeprVP3gYZc1+Fr/CnRdrcGA0DIu7CIhNURrcYjfn7Qr/m1cZSYpIs8U2EGB5Vd
XQ3j0hUgG7TXYEG1yUsQwtvfKJUo01dRVxXfUQN1krMiNnaSSpFSFtJBgF0LDJw8tyBwbNA8VSPw
3SVGffG/T/xSkhRqSmArn4Nu0Qg5HdbpYo1FVGn9I6U8hj9fP0RgJDfkSUZiqa3wMaFhbSI5zfkm
GaLNcBQR2XenoJZfDrhd9fMd+y0koOaeOtMw7i078dBD63JfQQupEmGMqqNnk1+UehGi8YTG2QK2
DwOM0qb4RkDSLW9moEaJxbXV4wXHbGNvuYs6CNzfWgQYb/V68qh+UDvDJjz0J8M5bpVDyiQjuq0e
ngWXM1TB842VZA6wZhCkNdgcaJQVYkGOd0JXXrXLYyONZ4UfO4DYjNPaZCdkLZwVoZxGsyXU1I7W
ZaXiorBb0d9KQCe3SWbgBt1EO92FbWJE1vzJqra4JL8uZ+QB98UGAKqLWx6J6qazuvKeKbolJo+J
Rmy60pn+OsYGtkdD3nP7zgp38cprZ+4ecW2ZkmQZ5Ajk4pD99CULhgmUex/7eu6tu8/Tc0gtouV1
Z29NNyqnK76WkEmm1J/xtZU0bK6vYBxjTi19DUSVaBYhgYABMbSBuj+8GUHq/2hgA8vCJvKrK8de
QaWh1DDQlf62pJaz9x2n2H96QnHjsxjQrtNCCVYX8L61t7NfaCPWseKNenzn6VQZYbemJl5Pwhhh
F5DAmspz1KYJ95tj0crdisi6sLeB372S4DZoXjRlbP3yctkBwZfmFmRYX7LLk1GcFCjFAJpoaGXH
+4Acb56vQSnSFnVjV81RJjX7nqkk+FCJr/XcsfCLCY4xrELphh3B0z+ISbPuNSxDrbpZRerhgKZh
pcmoelAUe6jwyF1TALi8RQbNMn1XDG57r4HmzfHJNvuz2dvGaNTgkNGBdE3K2ZXxdrLDrN5THXzp
02Z8zepb59gBiP1PqA1vMwhBSirSXD77JrOOvr7ErNodiY56n/L/UXt/OJZ7C/LkdlKvgRYweLKn
InbME9qmE1VLTE1iqpttsaq4nalRdO7OXnWaM1P5otd1eBeb+rp3rELzjqU9M0mcNtgEbhZiQsf7
zQLhkTTMw5X7DzYDHNey0GqG+yj2kJainoqgolsePmP8PcG9vP7YSXv3Xihp1XRJC4y1DEONYn6a
f7RctwFRTe5n/XJ0pgxfg0TuSOkcRdx0FYdPAia4QoZm8XG+wADxeDu5nd7T1xGcGT8YSq/xAVyP
6j7N5Ae+vaA8YNEA30+xTmmW3/ghu3tWrdPBxLgIQClLx7ifP2b3R+a6Eue+ps+Bce7mdQnpT0ij
HfmC3EqrpGoNXQ4AQUJYXjsj3jAc818CAftY/503SqpWsJ6cciRUjT5JXFx7SSFvB8wv3UxMszci
faLQp9dSLToHgzPjrk5vRsWan3oIXH/sOcaQzbOEflqxTb0Nb1jMomrSfwKfb9TstvnnWQvSTuVp
zW+/3ndoUwRkjKC9ZHb+/RolDL7d5YvYxma5ZPZFCfkzX7NKttYrkZ9a7ZKrLwQLQnLanYm+5VoR
7NYNv1dGMCwT6asPbLDU/OKe/tOyTyXHJIQUrtimpMNs/15chsSXHpR6g5cR/NO+tEqo1wqMs1Fd
NYxeq/z7OIsX58XTxiG5BiAelojDDu15EyL5MxEm7mmb0I+RifvA+VgE+SiGRkddCJlUBWGOdj5J
AaUSBBq+Cvf7Q4RuYzbpPwOBl4uyzitg+9bZ1oTz2WfS11vuQ0XA4+kRreJ3zzfmDgCBctKq3aWU
sJSyPkiG/18F9QIUbxAk8+qx01622hkvCPVOkIObeZz19Aa1LWxT5P38Yq0APuHRwheyT1lURFXX
6ibcIf2ln375LjRD928/bXxp4IsXBoILGp8QLtJmJwCwt2OdYS6a2YC69yjEq785aTUzFwyeoGrb
HDpJB6X3vTXeplIyQZGEy2rwvrd6TfFNdDlI1w4GandMIMWlZsDSxB8ASFqtHHWNpepLhjhtthOj
7e1LGxe30qfrN49+Lp98Ip6Wb254xYPyvbsS6PxGa/CertWqqfHPmrdc1tsA4PL02tS8sKM41beq
IBHLfhkaBEcCtei/bLgLu1/zJCZ3szys1wRXZmIpWle9908ckOVovK/ok2YJ15TcqO7gprj6N03Y
7xhg8Q26yKUTjNoBHwteb8wD7Flrw6TitVh+jEcN/B5NntPVawM6zfcGs6i7nMLCl2pr49d7rSnR
t9173ybs53XGYLPFa0uOKjKAbXpcOm/JZ8IcV/MvG7nYa7bqFfaRWlY14N3WOiE/JM3aJAXLfIrK
tskxNacZ8V4CwU+cO1NM8bcsUDnlaS0OvBtQPNwNHR9R/0P3jJEAygN5efiRyrfgzyO4SGAI07Ao
1hGdzbfbYB2mPQCw0rlvtIIGeYWYe/JH6wsoON2izi1O1E/6CxD+fp/g9XObMFQAgHQ7qwpwJBR3
hpNQEa+Y3Z3/2qpv5m7FW+louAUbn+VhQItnt0UgIl2CDD46xwI/ZIA1VPGUL26Rwc0Z3KIsBiio
+p6ixMNnoe55GiQ2wkHXm0ACLa5MzUgNxO/IQFmYBDzTThiSsbmQeEwxJbU1kwq7IycfMQeqf36o
YdI0F06lTZiJybTGNFi/O1vYBlaogbnKKUmLAExJQSSi+ep5VU3bQib7Vd80APfhhSadEMNINoX3
8uz/CgIGa+Eiass0VoBLpCAxJV0A1GbTpZWo/HjpsuDtM7ymQTWoCU3tYtEb3/P9s3ow5+Tyz546
zWYS4/R9HMd8w0SKrQcGUOJdBHgTry9eLQsTssawlw6CdQ1R9zlPme6AHU8rLuh4fItxL97qPWZn
N8NPVFsvQZgotYeOi7SZVrMMRhkLZuV7NpbWAC6CrVozSy5wa104VWPTx6hkT8KKdgHSEsKxbVeb
gnseCYl16FrfeanFkIdpjgdHdEIcO4b8X5RFM2WNRPUIOLQ4E8BnYf6TzcYb89JOi0RH/epgRgCw
BOmDZDC2olyrtq6VuZbxsfJ+jCeqQVR7NpGkHuqAp2vZ/wFf1LJ7jOVKkEPC8jbMlJnF5c1fK8An
JmRfiSOpKlp2G4mbOMnkgpXLS5uXI98y2/4cjXxf/5ZD8TyXWi5ABpNMd8XwaZO685d9UW4dohmB
DP9nF2uu7yqejoBrJtXubbSdsg+dZoiHP+8Fni7nb6PJZgm3Cs+HBBWU/CR/wWXT2TepFSQtLj3d
or3kq8iofL04+UFRqB7nYDa+0NXbvcDP9yk7Cepk4Sbprqowy1sbRsnJSv5GjlLc0KHoxJizyMZF
iOU0dwTbe9T7GSURgCiSY32fDNknBs6vraG4/vT9c0CA06nI/v4cPjcy8Z8yL75Z/E54u8Tk3uHB
wd654ILzt4c916mUTEAu7Z5Y3PSSFsYpvRHmF+KpJ4Md75qUC8aOZAkrwEY3OzdMxD58P9OhW5P+
otfv3EQVQTvV0X+o8W5B8Hm5wRUsbt4oo99/wr9l04Wvc7cxuvyYtOmy+gZRBI4bjNIEVA6aGRX1
qUbwgyKQAQOsX6Kx4WO83SLqSyxtcJvVKuvho1V8/H/gYMhKDrTVCehoz2m0djkz5DkDImnou4mv
Bq60hOm4eQTN5dS6wCIRJYrFyRu1IWzmAcb82gdA3V47dsIh8xUPDVLvHCkzqZuq0CwyjX0WRtAZ
+o1BY89ZH+t4wIgfSJLrGcXOHvt5qUw5+up+CWdFlw5oldmTXeKgqUrgnNGgd5/IGNec6+n+41ss
ayV0yG7V5/6evVcZYvLmgqAr4fkOsAohS1EeW0VSrtiJvANu/b0py0e9ra/m/6m9XW0X7aCa19cG
WVYjaxEHPh3pUNjFfJ+cpk8WBr72f0sicLdEa4XYKAJ9vS2eRrDFArRrhp/5NOI8T6Eq2e4SZhqC
KljZ1r+m8Vs65dN6x6tPvXAvv5CqkykSTPkkkse8rMFaxNbu49yZUpw0F2krhpErG1gdmuszrcoe
AlF3dtZlF2xDJCWcU3ZzbGkc4JS8RF6M0xrQQls0EFQIakRMPE4EUBzAMGH1sd8Y3aL3rLP8oeO3
G7ynAgF+oQs62GITgvxUOBAXpINdtSfHPjEP6LX15g1GpL58dx5iK6EaTy1S7a1q5iya50twvnQI
lRjh7dKbhTMEMESQpi1Wr1jE/80MiK5t0PMKJsMgs13MZgQTXjNzKRtZOAW/sTB38+cADWuNzU1F
z+LPcD5tV4yGJ4jyc1HDhbj25slyZ2GjG+IIplFDZz/WjXMY1FqUTbZy3usmgGpbWwDo9Vr0G1HM
nVmw2HvWqey1HrvhC7fw5fKFUXYWq3jbAX0Zb6SwWAS13gDOy1a0uvlO1ziR6hE/qnfEL76rOmFH
y1PAeA4ZOma8Sli7t+ek3BNVs4cv8ufHunqcGyKCCw7ExUDg62XuaTDpdbbIAoR2Lc9nPzeIM4lt
HkhVP0ehUV0nNSXlGtDFvRpJOkn4blsptOOayTgFv9427znA4PM0blBsCdS1jBpp9ejFGcPVL9JR
0yO7x4wWpkBA5iyJhBgv+JwCqstiuI4xdBSFYjlDuIE1JDiJsXRFYpZggJxSDVAZv6LSP90ePACh
c2IljKDx9lLJ7io8qr90fl/Bhi3dXTI0dx63IG7FtOClGvG7QUFWEMVW0YSQlYSJryM7DFonevAE
5CQ/D3XoifYUsDUSvoqHNHTq6SymRjOgBsfs2X4ESDMvz6MQACTgEGI9zmauVDF4QccayJjV5Dnq
yZoHA6/jma+Q6TPFDeh759zM+U5AuTAR+yyKiWvf/T+c/WikOo1bODEid0l5i4IiuzX/u1C0//aw
pMs9kTMPoBA7e4S15TcEVaaLIedAO2hu/nNvNAPMtQLm3EgE095iLsG6qbISgAgCLm+5Z4vTkiL0
gsgGp5TOTpU6FyboDSht2TwIitCDQtI01enNl1jX3mv1MEVxLQ428N8IlD9OMT8tpU03E/QMd1vX
KlrNeL7MCU2IoYHv593pNeo7tCp6zlqLGuR6iI5cImumDlI2IxGJKhQrZS2168gryLxcEgSoCTKK
IA4cun5/Z6M23M5Bmtm1Z7ja8iURgXXZEvHuGNlvGPQxyL3d8cSgUX7kJq8Fzmmo5/EVJPuekjru
OxJKB0mrMjH7qOgAql7WDgM7pDTrXJd7/nh9/QbWR32/IR4GJX/Sc7zpzBaFf8BV5N372icipQ2g
1Wu6R+lpvPv6zy+x2tix4QJ4TOX+NbtZsi+eWM0J1mFa06pHXr6Fxd3AppggVcFcNUjCY8u64yCW
AvwYomFNJKcJs8ucKbPz8xs5XB8y/DXWCh45qb0EZ+Dpcc9goLoBWtZW86xVRJqTZeCKQ2jWvc0K
v682kRkx2QfZ7BRvt+aLebMgkp6/pqcOMr58BO7doW+kbd++RB5D5DdftIcplKcqco0K9CyQ4WKN
HGovFi9cgvclqUXeJqb2QUxFVA7OVq/jmtCJ0KU+EWjs1o65iwFWN9s9Xiqidr7KCB9v7ikfWeVL
aTgngentsRQsgG6zbWKN6QhrPAVwxdTdEAq9FUOZxzJ5S92IhlYHIrI/Qg8bL6YMkw5WqoiuOd2F
Hla/ubU0STDK5v3GFlSbx30k+C7PArgZHkXvH+CjhAPFkBtl/F+l8+58nqlwECsex7xq1v9X82lS
bptRHfrl2XjpWYOKJiwW2BBnmwo80OAjTxpKOVHls6q0JLC/DaTcBWcYjLhykfT6zzZUoS1r9JSU
Nxgbny9m23VVrA+z1Een132VLKn/2XXx/Ad9woR/umNt/p93WrXlBNLTFHVJKUSswnNtFyWbKYPN
YWqEZLjPEdEkRhZ/XQUqqwNV57XqlSh1G047WPuqN84fa4TV4na4Fpu74hFp5zGehNWhDKVZ38te
ssdADPXuETl+fvVrCbYQHf9Y3vkxulGF+BZXz78sVQuJ11+aSHpVQtBozgTW8y5CW6XOZeaXpAmW
2xb0Eewy54Prt80l4tTe/rl1rIESLzmIFjlW7eb5xUAxc4Thv3UMBEaf96A0yP7hv0ZSsU742GFL
w3Xp/AdsCxBaOBB1VlcAphSdaN7PF279Bgcv/NySTQVSEIRPtauXlKRjzTDt3rmbZbPWAMW9bh8Q
NfdwiF9CRdEkDTua4wr/G9lJQnE70vvmtWhEY01dqXxaf6M+Vt8a7/vVHhtRSO4vYJNmSMNGAchX
85LPNj1JsuLsrIbEb8gLprbQd5S4d9Kdj+C6+ffOLI7V8V7dwVG9AV8M867CSk87gHDySFN7eC5W
pBrsAt12hCeUbtSG+xnvjO0DgGWnzpcgw+5QrAcpb9M4as6kDKdW8y5mettdVIW/zzyooXXaJemb
eXjH6SW3prh+Aj8FeV4F2uj1TzzwWJ4A4tiwXZd43qoonW89Z81wfZ3PZNsSB5jeJv0oWbNH0NmO
dCxA85t8zTTInsii0N/PHh6jVjl1OjqrJQRysrg85QPNVIDA19IDWfol80wbrAnla9YEwinxUtDb
KZVBrOBWA/hFOGMNQg+SpTnes3XvDaVChhQX2F2vtpSRoHXCAx4L2GRT+6UjxV0TfB5GY1n8kkhg
50H59ZOxOdwXuQgF3NZ2SJTvwtU+COgE74s0dDApXV37MDZyJINybjKNdN6cCmyijMTArI5cteMR
UEjgQjlaSvwmsg50yH/Np1KvO487okgpNegCoJynrs5R2pcy6dmqj02Cc7/XO617uNjk9i+JQIpo
vG/mSLaxNcQOEpeCwaLQ+Igzic61ki2wlLQlMgXzA8R7GYaZEl2SoQqS7r06ExoaOvcQzBPE8v1X
LInsIBKMWn1fck132ui7xXbmaoZrICaIDGBbYsJwV3Trzi519zrmGzTnRJF/4a5uiH6tH5SXWlio
RtpI+VsQdwSWBa4PRMQRxYj8A6erBzaaS+sGV37VtXy6WpHPCstXmvKy0T7CHvZNbmnrb3AGX3KF
OUXrY+uH5CKaEEi5DG3H0m+t0uJEDV3TWnzw69NURXCrNZYmMebleiRKvWgdH27dF1eMLWt3Ftew
bPMYkCtwdVDmWjK+Sg/Em1sHkY93B7Ft+aVSPvwAyHOv4jOemlXcNV3NR1Fp7nRmfdCysP+IGpnn
ULtGuHc+YYmZ2k/FXVuwNE0x1aUp6gk8fKclVwBgfvmgrkyVzFHRKaDRFhxDhp6OE51332blJ/wE
jR+4k3ywRENeVzgxX4GrfxKusgMz8qUXN2QYToXyHTviblMpIGwTBMepKoaxiKs0Pm4HcJ0f3S5Q
4G1qkBOAjAqb/YDKZEaiUg26Q/AaCZeYSXHCp442vpafJihWms0V/RNrKSmSKFOb8VIBPtLk0Qin
erBDjupyY7puf/T6P4k+MpnpBnOxUdmDLDXPLgVdL8WJHWgJ9t4o1UKMSZhtTCgtNhOW/gVWM+h7
5DWqg2sdInf1Rys++ljqUJrm5xLxsAfnPGYrVmuo7SfXOaKgPmghOmIW2433njoiMgh/yBURBxsh
EYemuFIAm+MUapS/p2buYkrB+6n3Lc+YDr6voLpAh8QHGl4NOzKoxFIWaUW7ObmlCM+R3iOYF38S
9SyOa0mTC6bpmVgG901tmjd9BiIEDDp685cF+OOTrNrGcENDfP/r6d6M1mKTyS/K/WslWIIgQsIH
Ujfjf+7cI7DD0X1cLwqJOqcv5GIAKycH6tT7SX0efKfpZaue4iD8bwjKckIciNcPReAOoc1DOTKn
/2SsWi47G95kKNYu3qaRGypkNF3K00ER2ic6hXapE5NfUs48WW9Wa+PgSSYzjpRtBAtJ7s+COJUx
wDizJI2OKvO5SuJEghpzzKWgaoEphxIrp0RTIeiWK50twBRMI45yGAt8XIKJWU0h0zJXusTnQf6I
3VrYvXH55o84O/aMsA3nfZjZctzkZQCHNmsWyGsvoIYyRD36mSFDdHenKJ7SG3iF13fMsRLwtf6z
J/s2OchVqifsAfKt6GMXKI6ZzSqnwTFp1qE4YZ2tQgilkyWZH4qTuRhGR/U+4gyi4AXphAf5J0Qo
AOk3ouV9Hd7GFJNRgsH/HjhPfoRjb7dtjI995zo/75jZ/uKwnY5ANBqCexgFjtGtqD6CLa/YhUrz
tFDtl0lcXL0bFi+w6audaZC9X/P2Ydiob/i2JPdvhjvXtAcD2XzYXd1HZJHW2hHrP4eiwfXdjouP
+3pHlG/9EJWrcQSFomIOBQs7y77I+UtBy4USiCH6+J9RupPPFdN/4PuAQ7kbTMnSQUg9Zo36HD0Y
qNiLVeR/deseTf3j17zEoKrQ40PigBELyjI5OOwUCGj0LkaxMAbH0d0INiP9lQ0scBGxSVUSpWhQ
hprWxuGKhSKNqbsNZVYaEGLFkLg9iOKPm6DH6ID9/ACudPtljrKYsGE+YLTshIlUtx+4qXD72ZoU
+WmM51TFYwP0U7n/KP/VhZUZGb7H0RHGeJOkaPPiUNGdTSDlfoo09cKXSFOlqfXU8vTpzel7gpEk
TKxHhmmMXAVJoDAmhpdktVsAUusUQCjaQZwHdZkhOS+4GT3PEXxbC2BK9wuPWvsaWAwc2UnRz2HA
zhUyoqoqVym1jdYQFwTCJBqW/jHBbui/u16bR8M+ogGnaYZJ1Ehnzqd44KIeFDc0AoR76QXwiaj7
zc3MBHz76LEp7761+o/w3y/WureiOKh6XhchM/J5nzmUuLq/yZjKtDBQ83T/3Y6XARFZSB/13vnU
+za24m+c+qxE6BQzWJGJpw8mnjrNCUGVbEgHA3d/SmX7c6mqxsfIoTcNGcoRbWeqrsJlm3cTjJ1A
wmfV+NrD4pnpa1Add181GBX7VuQCmTaf5RN6lzHxdu5SRAoqg55HT+sPeXSGfJ3PulfExNsgPVLD
RAM+CPQ21IfhBbPHTPrS40kgXWVYVx/0gC8yf2ffP7ZfHEKmGwKefvFBYk+5uKBY8ZWYTwQUgxJ/
qSXmRpDinTilIKgKYxA7BgRqY0QLcNBvsK952SUPDDxbTvzZBtV9rNPZVsDPfkbgggz75yK9XGG8
B7+CyjApxHiAI2Fq5y43StCv+D75rqsQuZTv6GmclcECl+L666sKoVcqmg3YC+ApkKRrg7OPs0m1
Pd1MdLNF1x4f6IWi9pedkDrcumU0uF1OQw1ATQI6QjE5oylrWJmi7Lxh+eL9xSd6atMeCo6Vknxn
x/rnjVLVCJXC93ufVwTbHnQhJHmJEAicVO3MyDFX+k49pJFZCro2DZ/SiqiK+Fn029Sn5BugkSgR
e+pdMbdYKLh2IeEqI6eGeS9tXS7Uwa6shjAAaVTjf6m3k4Pto5vTeOTpEmMvGsgfHUTELvBjfipy
c2gv/IUih2uetrtR2EkQygug1BJAP+VGNv7AXxBRD1WO31ZjokVrq8VhvtsCdHDw6Ygs2QYz6oZp
eOtBqr7VKemelLIHqH4n8oZxknTKLCugqwWPdhMS0gbSmKCA53m+AVXtefeTJUjEQMMpbwQxdYIy
R3K2XLWBvLrsYZfN885WiqXkdM844XEypsXUa5X8QM5w1PAY9GRrrwzHYoVKuCuYu7wH3oXO0fgH
GN4xvXDGwEYAZIZD/rcYe/mvJ7wu0XahZPPVCSwUrA27k6Cqks+1h7k478wdIWBF1vR/B+ODinQR
luIA11A1AtrwjIpHYV+hCva4CD9v5QNQUNgoY7VqwYSxebLEuhNhVmOrKEhg9FqxpkyaNOA2YI/b
LMPDsKVkfsfzjni+TIZAhf/LSFPAwNiyX5Ua58/akHGSpMn8pUPetJYX7CgGFLZEcR7QZMSTzw/X
c6otL3qoUp6lLusfPsJobmOWusTdp0plVB0hYOnCFnQgVLaND8SdD1USH2leydV6UAEufxqRAzTV
72gdkvZL2gzff5aEdqpys6/NwH/RMqsNaqd5hhGR+JxeOijopotPH+Ix8NGiWh+orL4WWg5S1BMI
fCoMNKSWd5ZdOkfg50jygR9ynjYtbGyg49p+oUQnNTsl03O5vGn48c2X0VSJrVe5QuUQ86u+AnuK
R1qu8wB0maG8OXDuK5WVeQC9/8VDDxnlK7cbpf5zbIWZUXRIVM6BNyF+kINbeNPVYTKhHGCziWb9
uDk2W2hKCc9EyLjaQM8hpT49XDmVs6y3k+MXjBbc4+d6edjO/5s12SWr6+eMVZLomY2qzhJo28En
9AdmJSrhhNi1ZdN3cspaYpTtV9BE9VUIc/1FJml9NUNlzfhR1FmoeD/+ozP1cNW/3YobSoSdO+FW
3lg+ZvKqWcMO93FRDT72KHMmKPqmyGdtvRTPb5Lg9RIfOoUziAD6Qu+FVUhjdP7+LDBSFWehGrrX
WR0FZYU2CcY8AH1p/pGbhlTapmA0bh8oH9cw0xzzMeVs7qAiz9Vln05Swo6oRRen8ddVENxHZazb
Zyx3vaec0TYpzyW5s60a/kkTm478s6sObiuyEEwLNRq8dpX5bWq/xUxnWLYuXk8pgag8avNQ7zA3
S7/Xvh4e8UGLgcGrV2KoVSugBGzSibC/Hkp4AQA77KIOZ4IHfm5n/rancQPg5X6r/c1EfoPkDKp9
wqCSxu/oB1EFnH/d3aOMvGdE8JLUuw4A9+C+0gbootglEA65pssV4oNVOWwDKpczISdFhPLeQhwT
nNgrxmUucaYbsamKlxCS6VjHAGq57neYBG3o+Bg+KXDd98dddTLOB9xcN85+OjRkyPThpl/6mOBr
jQ1veisVVTFsmsSffbH5WDdU0pKM16u5eCzs+xrP6zSYYYMIOsZS4dGrsR+f0LzkMzfTpjIk/R9A
lE8wYxqVI5XPtCMUiwVXaLzJBoq0PTGTDOzdAZvB8ndCisHlUC/dH3UlpPbAuM2Jfr+JhXGsZ7uP
xbur/soOYC0UlGXVjmRzffzWcujsuuWCnQLhCf/U/6IEWQSLR1ownNpqIMH7GkjopuZ5X4fn1wtk
+bZqEkwyToQNcUcZOe14wMDv2wbBHvqesj2+C3OM2ZX2oHYQzbd30tg/HOBh81yCaK0jxnaxnGto
EXSpO0PP2M26ghHFQBQnffkOtYY9Xgw0BJGkodhJtTm3XbbBayQsY9XeCSB6e1jOw8WxOKt8ot2E
SUXWeauE/wn24Zz348jV3wyZYdm3xiO2fhd8x6thgnT4XlFRg5Pw8kPCqTVFq1NtCr+3+Ezo6gVv
1eWagx/OSnLzCMti3cHFOOa5pw/5PGauU6ygJzNbbZmLY5TPf4OLp2V/VW/FizW+AyaSikXhmSlg
6R15DvmXbnZUxjaDD0558bWz1WA6jYrQQGWTxITGs8HecinEixIx62OHnNyqG3RFx8CYUQttvkf9
y7XejMnSlLwipF1gHLKfYzoeeD2P7pDHHdKDnMttmnjtOrU/ZFfjA0yT17oiYwTIjpNUVvlciqk9
F807+KYxJW5Co9P0NVGWws2eTSqwgcvDLyAMCyXPkbRas7dfcUGequi1m1AEAyO5N08mPMU40+4H
zNebynt11T9LdsRhdW7+XeUdEG0f4VzFMF+O75tUZiKM10ExMTMoOjABUFLAdgyOex8KIVvSYg3n
H7PYBuOno/vAaiW1VpJ3V+eBPKu08+n1RFKwpOtBPcrD22hEZ0wuMEuoEY0W38tiSPK5tOzhzEH3
lHPu02lVEo42522XTALwPKzeuIUmR8b/DpWfGPQ2+HewbzqdlwnVNqM2ThmtdOOBwcS2Xzlx0omC
s9Z7cRivZFGPr32Mk7BYskL81U/1r76GOckk/68WtwmHmQOmBJs+y/pUWmGVA64XuBtjhP7oogTw
r4KvoVRoHfkLlkjLpZ7sGfMaXAtU1hMYUfbu73IRpd1tEP+FQQyNUs0YbTJRYzQIEeBtJ/XqJEHB
mjOYh+dxUF42eMM04b8bwxu/uF4hwmMt+KX4w6pnpv5Y5Wg6JpRxo/5Gr/MU0U2Mq+denBpvfdgm
3T+of/UPp1/OCZVNxk8Qk9wYW175iUHS7Z111Hkl3A8QIjbKGZuL/KqtsqUH7zZB0b45M0gTBggf
efd0St35VhojQQ/WDI2nNyySZLAWmxJHle9QAkBRr9e2maeBX5BCKU6vJhaqYocpVloi3BEDubxz
tYmAcYcm7fAvhuC0f9qw0Pw2VGCUDSniBZ8HM0kWaLJXmGjyN8dS7RWwXeQ7V0NLu73enMDr6x5/
isl5ZBoGrBtwf1iABRISK1Mrqw/EMqUAwgDniiosZYBU1j7MP4xdyFolvP6aFnHuhVKTiWarT+Ao
11vIjqm3iO6bOWYMCjrp9+Kn+JCbCYNb2UNc2eDrVJowmarP685eD2F+VSkQn+4gB6HFjP6kYkQA
eUj0qvoPzHJA6ylOrT+aJ+PHYLUSutlsxO9Vjrm9XUaVtT5oX/g+WPobCzdKkVlqBHnrgauKO1sq
r9Mkd/QKD5M33VtOBehvWw2NiqYuEos1fyUHEjywJLocxZrkcuvEn0m6mlqHQG3avANnjsmObCsV
SwQ+NAI0GmwvawSNnGU4H3joTRxOvumH8p61QiExU77aD2vy9Kz66nIyGxlXQsadooApdUne/A3m
wKuFSS5ogksooziBUvftNiEYYAMCpWgGIPvPa9Sbex111vqX55ypTAv1UDTUpi4O/LlU01zHbext
7JPyKQ03xonEWHAt8YIVGQewxUlJUt3KOXf1YcSA8b4jIiLyImuCUjbaXxJ55AMcoFZk0/hs5Nd5
qXbbMz8qHRmhwV1QHy6AoyT1Tz8IXiLMrVKwLt2IjvsvHDaO+NNt1xp3tFMU7Y82N4Gsb4H6wPj5
vEvxAp2ECFciV4b8+mf0z7UCWXSqCbIhqX2BPXjNQkiKYxuY28hTFpVFrLcz1KD7IY878E5fMB4R
6Vr9xafZN9fO2j3cELsVLSlaDauxWYGFxCFPnTClWD3wxm0DImxXrsk7Izfd3uJKaeoN+zUAQEwg
IAnAlnjgkXGtXRjxI/MF/QoTbbEmMYeNUVKNeXgxF5kTCs4A8KmbbrQMO+2eWS6+ECbTE75Rjy3r
f7jlXxGtW6t/rGpAoZVnDBFo6AS6qr0GgpwNnyrG0g+lwkOguh+PizmlB+8gdYGfVQSQOlJXez7t
i0KF786mh3QALbLaOp02kSFLBqlbOiVywqNGq3SunJZKrJguteZrQ05hiQSF+qmwvEIxyOOmmeL3
2R7OfSkf1bWPojVeIHDmPymYAGWbWqgF7e8qPGIQqp8kBiqow5LzbLfaXu91AXbTyAq1/SS0p4sH
2Zy47SqRaDHEaoB0uypRI0O0gZUmMhJ2Js9rAJdpPcRyx5hWWlRZ9PT7gWsXNIRZPI1CMrXWkgBm
SkJ8w+7a7WfwuJ0Kz/JbdKIeu9dZ4p06dkGV4LlaIGJ0Ki1dVjUvelKQBK7W9jVyrLPslttI5iAD
67g/6yFOh12pu6EopjPtSv4KlowntZ4asercJZb9kUuSnxxMYQDlKK8QHWIuRxI4++zwfYiAMzRz
yczA6Xmr68J/JH74HJAsz81SbZ14I1dm1X6fdgn0uvWQBJXx1Gcb86XQpqzD+L/2lyrsh4bgUkqA
4BLPONZEcPMOqwquHsAvAaaRiQu4YpzcnOfFA5WB091X018jdoUaie28OOhJ6HDIz4c2jys+fc3+
qLuS+8Y3RJ5x/I3kSWZxbE+2VTVM1EWrmaFhNOeLG7p/8OlGERsP1jbxpSceBj6HKSZEmz7ZfVtE
ao4aNRSyYShEFWPedh3YaSZuC/Go6ODqFqC2/JXEf8OSQL/KR1rGyz+IC2tafCsxhTZpAmYfRDq/
S/eDD+An+R93F0DOhincn47loxZTzYdBf5wH0A0nf18CGJHDoedCW8XgGAJ5UswPMGcvHQEWHJq0
Yhd7NAFH2iAilB5Jd0M/vwjYFSTX3wBPxqyF1Tfp4fNEsfiDIAUmi5hyyIhwLpQB1t9fxAezuyVJ
3g8XgyNCxMAi0GV4TlXcu9tnx3LpViNf5byWgjdOjvbLksQzzcE7Gg0AD1ZkWI1BHaV7b4KUbMKj
hcURIDuWK8N5KUdxJXFZYGNrLUXEShq2fQq4unR1q6IeHVDJCgU+Wg7erDxb4hC9x9EbD0Cy1N7/
cU/Nn8T4Mo9ISsLeWFAV7iDlYXSjnMvyAWRhASkeHV+0XH8t/brN/9lAKOXgq9yf5ai3Xr2EFCjh
g+ZE1DJ5oYSnUjUojnVfgns24UIXOlDTdCz2/XXujrH8VKn3IyLqoLLhQO5Aeqm84FfHtb6uoMcq
PgX0MnVH3bc/y2tXMimQwS9lcVZ1Dd8rLeXQGw0f+LvXPkdk+TQDJDL5GhbWG9NbU5NVUnppHjUv
JLcGOqJ3ilRQ17vB8hSvrEiLjYlacsMmxqbcQT5+VNGF7ulw0gQjZk/AyLwa2nizf1ZqzBp1gH7g
5ZvBNiy2SHQvZJ4SxNP2jDidxYSBe90BqKg2hhNu3lrilyQwbvYBOEAtM8ntRX28jhOZNwYge/el
ZKcTGbR2SDs+K/c6P/Lzif/NS2N/YMAp8vFlN0JJnyf3E8una55qFvmqXKpLR/dl9gMIAc7ho+14
DWQ4uN33FlDLruxyfLjWM86k2BuSDMKq1m3HafNUmCCcnUaEYgh2Cdx1Q9JKE6DniTgMdpyzVb4s
sW6f42UighX4g/Iflska9RfpUVcBoa0znEiaQ39NJKOi1ezJ6XMHXSXtMuvS3g8A7RwMfRCOMlU/
zx6qIy3LZd4AxxJNcXwVFgoLfSTBSQLEqGOokErOqobcl8klDspwqtnnRqwE0hT5tvM/2trgxwwx
BM4iQXrkJSshLvh0wdRDTS5Jg2sXQXjOwbthJ+P+zshjoOiSKSGTohiss0eFv9i4QUn71mnXQ3d4
tQ+vIz66pcdQIgiGilgTFjRZRNl87cKuwPPvf29UO/zmHf19H4myWdk96zdEfQr/zBc4/iseZU/n
o+kHzstijX++gN357vxLavgulv9wfsqMgIMn8Hrk7XiSh0PoK0XmpiM5CIo3AjP59w7ePGcY4NaM
crQ+M89ckGmU2eN+f4dzpS6y3cvdgc6rLDr80/ONtDtWEMEj1dE82JIuOLOSKEXFOV6BjHd/DN/R
gbW2aPGo/c4m+0crJ3l4SBb34Hh/qOVaI50PWpGOp70Y07g7IdFp733mSNSrxBRNTP1M6bumfHcA
mwqXu6lRG/HR76C1Jws5c7DYAQv0alWQ2MFPXB/Lx5zBFvsXGYsXH7LdoHSXFW9JrkhypWkbpGCF
ia8fOP5qq+m57LGLy1HSNNkmf6f5nOzlDN/dPmejTJco55N9QPqe8Cc8k9bTB1OB1OjNnKF/d7zw
DGpfl0VVleaU5vUCCCgyltceYnKzt8pQEJopb9C5y9ZEp4/0IqIBGQEMBJFf/s6dMYWuMh7taLDP
Snam79HWLWeOQzj1CrCs5EAuYQIebsSlJj1vQdKCo8L90HBq20o+9uUpVRNwnmZPRSW2xKHyzBlR
rHwQfl/8wZj0dBUTgm+wM5t9MUEwN+KJCKhRHuSd6dHs6weBfPMnGPEXbLknodQWkbHNMBEYyB5A
AYxEfcZ5XqrKZuO+lqSMbjKaCX7B5+03VTlwA2D6JqBjvSmN464O7TDwNdhl6psqW8/Zd8M7OyIA
+OrlgPNuFe08t+5YMTxC+j9lqhwEsCp9qGSYlzfGqlpZeoQ87B5wfxb3Toju0yo3TQwYag6yjvRV
9Pu93REqoulfQQaLYEOew4GJxyeSzhrKY3SV5wGzK8gBEsKmxXkvohj5lLOUrYi2/jYYZZoJnkC+
HBKUtQqA1dMuLMcCx9/tKyDcCW588lrB2QZZYqNzGDnOcJAOgRhOnnMtv6qmzg5HVIwwvKmh7aYL
n6GvihVm+fcB/lRpOjOv/jEmKzHabsjYUeTyo2BH8dQQLoM0TsfpJtQblXXV1f8SQv3ZlVBMrPkY
CvM/jNncsUZQ8HbGY9G0enzIjdyhiTKKmgk9bCpi1ZB2Q8dyNgt4l0jc7/+wJz6WOM5FMsqbHcQv
SYbJVRQhk23DIeOCn2m66XyPibozAbslR9WXrnIblStbpkEsDrPsQLI3JHgEZMR1uFxYtrFdyG6E
ijLbBPTpFvN8awZjYrvXjcy/Ko871XXNvXDOAosfBd+z37T6gKI2EF/W6+L9KrsWE8P8Zs61jzwH
fERKqTrlKLKlTOpx/41p7Om4xA7UoIbpL1fIEORdIOs4+cSAtH4uKsZD4Hij/V/BQ9HwZBgmxGM5
wTAAN7geCtESsHiUbpPyiThOEub6g+wOY4J7XupOxlcFdKGvtO4RCRY04E0neSuHGXXZZgjHklKh
cWssVHs0d87AHoWf1smr1tcq16NkBIMX2umBR3dJax4KkqsVvKjB6OxrwiaE7kjpbfWJDu10WNkz
4zpNWnpbR70dxZ7DLK/5imrr1m4PXs/PnI1j0tJEUzgIDJCyv9tRi36bVPg/8xlW8AI1n/7MlT5z
z/rjDadkzHb+/+Tx+Ydz8TTcQtNPvMHzNXfPqqWhK6mRkMzkU8JnXnTGmiqaemntSt6m0TlGUfIN
H08tPxeEuIitDE/rN1ErstjD0B/l7hv+2PyCRJH1DBA6eh+PeOaYBWVkQWCXM59G6sDm0xSU0m85
Zl/+yJTvVWBV3NkGPfkpdBojATNFLnox4UWYnWllneVaYahGE5Iqg2f79vjARVKxa0+c1Hz5NWja
2bM5u4NvxtTQVbLbzcWdZUjXgcc1gl0hpIQ9qKsJFDdF3TbfMyX6JW6rFU/2MzFEMErumSCO8Ww+
C35Vbwfi8QylKhDWHxcsVr91Qh3aQiDXJAuzmqTTHcj+Hz5AyFX1ANHbFL0hOr7cey6aDEnYAeFK
wpkrlqH+JY119U1DfoZcjDnWlAiOs+YBodsABFqz/8YOlKxA8ofmfp1M4aZasn6a1TyakEqN7Fe4
cYFis4hl0vYW/QDM5x1yKO+3m76N3MQDZLYYqkkpU3sej1xANgMrmAkJuyvgQRzJdVy3ST+k4NK/
7SyQyDFkeVHU5bYlnCLHl3UGHobEYize1PkI/zWvjGJfX/luX/6paAXRLTkPr/qf+Cfybb9psiM/
Qq5CMWtY/Xk/PTQNWA5yfrUNbD/eBOsob//9VwHpmkVET0Oyn66aMJK22sWs1yBMbUv5OJhndm0M
BMfntSx1upNX9ZZ2sopqnKOeQtmks1MmcoeZ9NE4Mwhrx/KmGfDwE9S1LzMx2s/qpTcNJEyWRB/r
p9TlK0D5vMbzBX5bdpnaq6y5tc3X+JeduAP+Rk6eTl92vm572snpGkpDMIqUwVc8cYKHaWgxkTUK
r3oVnN4cDCqubfCgzwBGpXbATsrCc56wC9KUQYp+ncl1NGpR8x2egvx58ugDKvAi/8YITfuHl504
MBFxKs9n+PITdbSFw0D3HHEJndBNf0Hi/1orHMvis7O6huFn3RH9o1RYKHkCaBxy1xg6mwsUzECv
YViYVlUEDUA+Z5/APV99tGae6ZuDJgrMceeMS3flYmrPvcZs0kOIoyjiD24OtbsRB+UkpIZY5y0+
zH+G6WJqFl//yXkX5E1LbWotqzXrNQKIxtql+gkBxwanscK+uE2UUipSdJTe+v3P9tVZb/aXnjt/
4snBQFqJrOAYS5b7cC44PgG91wWLPu+Ts8j5NOmvAztyrWvUCqvX6cJlB2YPy8+P3UQs4HnnD5Eg
ywhPQDHtquzb0+LJFkB0VoqJn3QmdY5a50WdID9ABVYOSvQF1k2SL8W2QthfBOC1sawzioOswvcK
yhl3h51ybNOyjmgHWB0Qck+sVsgZJs7JLVKDTrJVpxPTnZnRbQsXviRK7R4efsCDRn9+ekbxibO8
RWi8ZnwtCBFHCl1uOtMhJBFKsG9UoNtmPcxo2TOqSqweEmX1sXnBI6VyIOliCOtK9gIMQNcDPWsg
G/ukJQJqSNp0WypqLO0ojsi4nk9QxY5balMMfT/QObKS7wueWnsX1GX5vcKuNDxehHS3A/0acAok
zamBrVwrKMnqEz1XiYYCqt3Z/zBWML8rkKa38V4Z23QEoYs3jXXzBZTVma3ocC2HRJ3PowcXaspF
WWiB7b4SlvKEe4VeIHVqTseTSsh1EdNpmWh566NJwz8On7kgCBMO6432Dq8yo2fc0EBtKI8H62hv
yDxNT4YYZfoWvOy8ioqa2LXVr5lrDWCq1BE5UNn4fj3rP/ecb0lLLmnauzwCu8uid1Ej5bpSiwUO
HY4OHrSTuVytE77WbR3NGLTOd1TWPjWGxREws9J0nwj1u+O4Hm7cI0ZfNU+MOc2uDVa0FUblETFR
QYD7DuTNrhZb5SrEKCyumdRuaYhuG8SAdqUoLBJWkMVJNHTqNwvL+axRVSBtUa747QZW+g7323QH
ZFxCuE6svxIeUAHbfiFPAFSXNSEmB+ov16FYc79W5y3LSXoBi6zJI8PdfVsIxGc+gnzlCvUag3HP
U9/vE6BnpdfVBSzC/2woKsiFXzYpRczGM1MPf67BxnH+9UuP3dj+KmfETuIFWIdPaJufXteBRnDE
KGzgit7pNwtjr0qRTUlQbY7vnbHzFQqCyTb3w+Lg2jzEI8bNkD61yi7tQBsAGIi3lXsGsOmqYfZu
c4y9oB1jnw5//JScns7U9SlHojnscCOQ1Ij4YI2aoKpCG00E3fTRF9nqwrctg+Va6p4W9M9ADdk8
lbkOv7BJuEl66sAyc46j5mfitmM5I6FHBvL3YbQ9c18ltR+v+1Kb7tJHiuoX8fqV0HjLKz79lhYv
BRMphhfkMs6WgXl8OqTR/2xTIWWdyVJhTAITAsQTeX+vHsWU8WcdZcElCDKxy8Okq86eMvcnsi9W
T+3g3jdu3zzp7nhLjvpOSiRbX3pNvgxepJ4Eco7HKu9WNoTAv0YLwxNKFPW55JXPPRwQvI/hOsfq
vqhx3gJqrkBI0mij9t8NcQE11iADVTNi4gZBlHR73p28+BA/tWHP89TfHZQftQqEhmPEVWSSQrwa
qBTDYGjJ3fvfDBI2ux4mf76IhIZ03fTxFcnP4v+U/VXDeZThaGsiazC1PFnRCL1sTp5OC1iATE3j
0tfDcx1R7oE1Sp3KhroLYsZU7Y/hGil0v9QhPPKdUSLimlF/e91GcxLrDjht9KNKvmKimcpQn/94
VcUNlCOcwr2WxTHWPpc34sz4N2COuyKpnYYAWStIpgOBe4NilzLtVvVTx08BxZ9Glo3CkH6CB6tW
nvMat9Ls6Qlz5OU6BPIneH4PrtQ7gaxKP0p7ei67rpbGiYJWJw/P0IyWcHDAeQ20dR1OugIibBWk
OQJNQvkqyH2VqAQC/FItD8K4TovFkCGUUji+lkASTp8bdiOxbrybu9mGv+4f8yXvuxk+sNzmJ/YR
QJV4ngidNSzGoofLFVuxKYj1Dce4Tg7iuHWcec8xVEdW5g8ZA/WpRcevfiVMPyl9jBcL6D32Ci46
bx6nantc/9MkN2OmXuEoH6OvUss5/Vcw01JNg3mogcU96O6r3plArVecioGys6T/SUh545KGMQLU
uZHDfZRL+Is15WdL2Veg7gm/m4R9TXX99tuCu/HYBXDBoeGw7DQZPJ7jJnu233ASCkCzT3R9e6xm
a4B4UiEx8VNl5izppDKnNmuGuJmcNZUkHnDLhV72AhDY2Qx7LjNioN1vFEJUGVINgOC+HeQO48Xn
F+C6qaC7yasFhaBtygnKq++Fiy2qD/AiwdIp3ulW8klqpXNeB2mHYpwwrFQwvf2dK0tj0OrtRvXG
9tnv00TAmuJDdI1PXzWfMYQ5QsD8sWhBxwqGezgtpzQ0q8v8loQ3Xe+iIpyuYoQsc9cBrQJ4eCfU
71x8fvuXbsk8zHh1/MPNaVID08PFB80N2cAw4q9MQESmxcV0iUOiFtpsKnMo9ZFyPh2Ad8Q7Ksh3
PtYjTGXEh2RN0+P9SsJw0oDflpGMtnleXxJMNbF6QMr27xU/UUR/tzt20drD1lL1NAT2PMyAb+Lp
GIkxnGZA9rEH4NpBfO40KuxWQc7E8vQdvtHi1M+mm/0TvLyuMjpHSHSBBdwJPYM/7JSrZ9ZFaHFH
AqYAAoa1yBVhiYsaIQnOKFtqg4Qa2zQjPX11TbNO8lEpJYpHEaLcIeZuYP1pL1X/J/MST/uj5wE+
L8WVvH+WOcR89d42gx3h5sK5BjRFqQrsBrijDkLAXXnfjUoOs1Nx/8kLmC8J+AHLPl29Tbq1KEKD
TPSTlBUPJ5WkmcQAQ3klOpj+gGSs3jJRHGMK8lhni6kbTD2qdXX+vZAQvGnFEZ+wZKNZUx4njouo
HT0gGALgqjIIQwqsmgshal4rxClTtue7LxiCAanMJw8pGUS/FDeVSI10Ka1W2BfP5kRfIFKl5GYK
3yundGARfnOdDGQYezodcohv13K7keZFqZ61JdfpDZ8kwti9Rt0FBv4l2u72VobzglCVsHf3yXqD
9ilQZa/dob8h0vBKO7lYrfcuasw4yNLi9HJ68L78CDimj38FSKeUpZgNdZzH648b3nLrkIN0F1wM
RP35v7k077KzS51UhArIHHauyn/yCUbFVE34JjDT9AnFNw/nxOIOikB11jHysNEzgXpgqKJ/gTpO
KdktJAPNsDnwagX+Pr2umO17DWQOKJnoggGXQEsaPoVFIqlq3ignpk8K4D5pZCZxfXyTZQIjX+T7
owj6p8zNhCQ1loXfmhMpD4+sPiKBXvpVbzJ1zsS9nYyMZziK4JRRxCn8ohPiGEVeLW8R78jPuN1R
aeEXrjcUG9qhed2EjL5x8U9n35MdC8rH4BhbIB9brHfgnfMLWa3cgNssgvWsvvVBdwK5Jnt47cse
RYquMPnMz1BYwOthylXssStakIaFhrt95jrWHGWxcMR3jb+I6mDnC/vYl7RI6+TgJOfN8rSNOGIl
s4PqfumWaymJoxmi7uO8OfRNh/SADWY1IHALCE7OhmY30TpaiAXHjjfd6fdle0cyeRlL8bwfGj+D
jhCfdwNgeAjEQTRC1Yf8UgkwgGkV6EWNOaULXAzK2l0dEqJauFPGtY3KwIUFi+V9ZObNzYbAMLhg
JmAk4R9RWbgcpjMN8uKN9aFVOlFc3MIP8JvrWqm67EYUmFYcVaIb1+BUlGnnfYTnRq8OwsOPMH4E
teUSFhsoavvUGgYsFu9T9LXvM14da0uIqd/ktn/k/17+exLjO+b0YUkdcyABRy9Vefk5UFgpZFxj
qrfVLInhs2gMmG0rez9JW83+nK5tP1mx/rl2M0HmTSCZ4hqMm/gqxKMnd44mL54TLGF+ZqisxPE8
guJY6BIXm4PuUXmp0j9EGmZ2XTaE4+orUQ9FXtVQRoWn9Jxq4jM0/e6vP1a+c3XxgaJrV3mn+qjp
UhMQb0w1MojVDtvonYBv10WYFKbazBiMvw5N0T+AQWRGbe3fsg95W3zsJ721NvTkPXN99cvCajWL
HnoJoQSCkugfsbRiFsI1+2Nyf4dLfoNxJfltDQbE8/+K9LPu4vNB6ylRK/qwqIIjt9Zg6f6Tu/tt
Hvsycp7DUUyveXgzpQNCoefIiR3VhPw/XbSR0aArHLaYiuL3GYgLi0s8wUftwpxS6/7OedE3z0PB
DHFaq6+mbBHHhAhQGBEaG40iy/85jzJKhe2MR6+9aGacElqlXJLk8+mjvLP4NUdhZNW8Zxh5z5hc
PWgQm2qUs4GzTE+1exP8O5B21JGYKY8OhfZXfBx58m+3KuUGMc01Kw4rlDTvaghlNW2j0yftRaqh
oFZVPE9w1szwnT8uWT3lxP3LcqtzeidjKLA3/XXzu/j8rgAN6RQkQlJiaF3aEQ2mMkYacLYPtjDW
c3323JnKvLzWJTs53DfF8Gdc3T+Hyb1b7opTSRvQkn+2l7Dny7VnyfAYvvFhJ5dDzF8vJN2mozXL
G75noiLj4y9sXXZSrIx+Pc2q48r+RJYDgd5YN9pcTpyD+/oZdJCRYs8cAWJTUJUKAowJvhAyb8j8
WMRrHMsi6RAQ2jM6psIG2inGSF4gh58NmHOiZAvjZ7xeAnYyce7lDSs5oPk1gn9iwKjli6kXTqtk
qdZDKTzKsr1VOQSU8WEX0QKaPCZ07Bjlo6DcNOCKx2fCFJKqTMrtGNrEU4ex9bVgrgvm5xCuFgkw
rtQDLGVPvr0kWItoHb07URtPYyFTcAI9DzIoJNQ3G7pH4Mwx788JNFxo2HqTwZ8M5bmoa/Ytwnn/
4RyhRK/gDF/tYTlbxDIDEakkX0gAhmEC1844nr7fanC004g+gpa92vWnnBSs9kQNpX8J3VO/n3cE
41jvniFXoKmOeznmr5vks4mjBgjq7nrvprFh0xB9bGORh9wdoZr5/8C/ZRV0GAeJGzCZ8+enV4Oe
BeMAmgRKejGffWkY0sX1OwBNP0BiNu/4tCwYTVtI3JGHvpjP8iguloUc5j6/yomV3EhW9Xt0K5Yy
+A/oFw8Mjbibfsq6hYQB6FpM7LCVVh9brBzKAzyjOpC4XfBcXYhGqC4wEmb5MPRNnheh4XhY22gz
Ki+IXdURchp4fvtnG3lF4Geiy4jsEBrj+V1H1bVBwM60ZhqTToLscV/G36nbWlLyI+XGWFXypOww
TofijJPM5Z65WVTlBaXPGX+qw3FjbWnw1sB0HKHFOIDda0EnUvjHcgO+o8BSsq1cImcGFd/JkaVp
A8gOeiM3xecHyL47/UOBDpf7SXXlmVhSukOV6e0j7IVuQ7kKE8mbzPZAuX4Fpcgy1niTjv++CuSu
mK/rIlYk9NFkRdKfw0IY4TU/SgEhSJe6MlW0Uux/tQptblpPG9mvwXe+QQOguMCeJSIWPSzmcRC4
2pBSfk6jU8yzBwPwRZj/DfIjvlFRU8xslMcwadYNqZqLBfdYuxNVssdb/nvIkiMX3LgfJaehki4Z
0nEK+yZg4o14SttMMxVfzZsqd0hv/WdGBWSirVlb0ocwZANfWAs1ZCzuGKyLQvBGYRvyoa60syj0
r/hMYUBSH3BLsqhl2g/qEuA8Hp54fwL0FDjgAFSptL/H9UKXjc+Lc/+xl0gHy78ZY9udJzZKvhvr
Y04WsDe+6i/T8Mt8QGIN2gKD42LoRfiaWp2SupYrmTMHKJ8q0Ze9WBouQt9hI1oJH0yjm/B02qC/
T2Fc01dzlCbpz6Z/RgrXHXVvbJa/lcR/1FPcFBu5lnWyDhkbNZmz8UZ6oNJkMXUDz7okWz2GwQeN
9ep9F6wkbUDthv/zGEVqb3lepeYGOBZPv+KrpDRFrBsO0RuvSBaU9wu8U1pmvutNByQXVCK7Q3S+
0d+fpx4lsEjSLAqC/6Gj95CYmBJa0ge+X4Xe3JcmGeRnulzEsuSq0la7E7DjZl15CdA6Or4beqJB
74ouMash2Gr8VccMohh/+7YpTS+Q2hU5NMNxEHCBfl1kFJWZpUPHNYzAC2WJTLvDeBqxinRl0SOZ
Wc/Iq+FA/qUlO4klbcKu2Qu1QIVovWokSnB7H2AmraGOVZGgHb0dJSZma4taP0FZP4GnO9g+aKc1
fkhrVwlNlSQkz7BFp3cDjAa/qwHoClYTyY67G2bwBsR3S3xRncbsQFiUl4aBW2wzp8u0Kr762nT3
ALRq5fwrk/bpQ2I6R7xAJ0vZ7Uva5d0D8sF4GfZ/peupgTB9BCKPX3fP4/40wRHN3El9N5XH8OaN
4kTM+frQJ/iS0VdNB1pKGyO3bb/5Xi9021Y4G0SH3B2SRGWtwyOhOTP0e1LVMrmsOsgwSgV2+x4T
eCnaiWppWqWQGgXNs6B2tLZjVITIxtfGoMV7PgxAaB/YiLEP0zZhkMvsGI67dehdTLgwkCQaire7
ySV4hyXbzQCNdZjyu6N6h3o6e36ri/4upqmVqEB5c0j6BaxIZaInFT8ikVzHHsTfUceSd7EKiH1I
DywANHX7nb4a3/nFz6L5PsvfKix7M0LxlBZxyMH6qZJv7sHGwnBB41unXZ3A2q4s0k0EoGsmnxms
R+GKhCzE7Bf9PSqJRGQ1CwTBat8dSZ5n+XyaW7nP/CP0IjHeHkra4IYg2zrMqjBgaQ7MC4IW7DNa
fjBw/8BMCytFJrtWtqZbOp2L/q9gnr2OBGMi+ksG+jZx2GAdVdo98zB9S/ACj3eetYqjqdjYTDRp
aUnzmsFykjhXBXiylLdgI1YNVl2QWuggqy3RujMCaZCMduNWnMlaSpirbSzeP9J4pW6eXi/coX2F
GmKL5YDqcG8SSJoPhCS22V+pDRnuaS3QCFUOGRWIy7uWtTaKmARmt4KiiwCLLXwdQF5vlNh2iM4P
k6RuSHlN4N5Li8BKPc9w1wH2CIc8BJEpA218jU0vLRXy4tssVuiYzKD/dBNq0vAJ/z1ZVD5HEKSF
P65BtqfqgiOVnUxSA9KVoTLafA4ubYFf9GxXqp5PbQxGeeK4wVLbfCFyRxRlMereJg6kx7a2229h
aEN+9i9B8C4VjMgnq3Szp8PUJzkqIIKNQHQ+D8Vy6fdYZ6i4J0lJlcVIMAcHuQgF3dFQXAZx5QRy
RuXCb2PrS0d5I9KDT3H6BN5k5hAjFQGAEq2uG1LxuXv660x+tdNh5xhXoG/AudHGIoawr5CtDks7
QqexCAo/DghhrzZ2kWkSBxd1HMCLO+P4DUysViywhMxfgixOqzhMhVRTy3f0tdbwoisaYbeA0B2G
FPIAMU0Ege6MHoaRQ4tvEaa6+9bqcDc2qn8/dkQIAN8QonvxO1flYvjIUM6vbjyMBh9wAoFaYXLE
0g3uvq1AXTQTq502ukfzYs4zSPnQhxelEJhg7ZrEELVr4XzaQNyojGE+ryVqKw3N8dvj1dgi/Skx
6Iw6DW8ZsXS7QEdKJNSbuaOra6uC3IncYWyzxeJmCgNtKw5nGTB7uG2qJLh8HDe1MtFDVAqp3W05
bzSd9RcgwvbHYqdT07b0ajkisEc/qh4ujFGl5rEv/1nJVpnXYtoObDaaWcpGASx6d/HRVlgjJQ19
CW/LCOUPrV2ooVaokfLZbwfmPG6hyWO0cK7wOloLS9EoDCZHMVFyrGnOiRyx+N08/yeAF9+FscTe
o74Mtuf56gSqYBTgyi463QDALV6VNsUyEcTNmRnCnv3l2Y7oAjJ0dj4Qi2DsdKusy+HhLwj6lqHK
XOMQpc61YRfxW9//v1ZF14/aAx7K5y6/Q/jDMJqUQaB1a/fqbHwhgs+Tm5TlfuecXU3zdqGutz0h
ZuzsUIchxY58ec1dW8wmHCbvj3KGeKLA78aLeVjwvlaafj6OXkwnPzDAxmlIgzTaUPTanv1p/NOr
nzVo4fJI5eNo6XIb58ocG+T8ik2hNMimRkp5fHjCnDfDINJhGAb/41pcxEvESvVkhUqk0ZwzGJbS
jTyJYHiRm89Zf9jBlNCK6fOIOHP1+ZGFFSohKF0BhZ6xk7xi2fa/ZJKUxIAbP+KY6/DfDlPraRsP
l3cM0hyBqxvgxmbiBEX4xeBNzl5L15rvGHJd04QgTf1wXPbx5uLHHNi2BTCEkmLd8draE6hpl8FK
4S7NJFMsiKx8j0G5xBGsukPoqDUzwDcsyprxbU4l+eQ+Zqz9KMWVqt65my01NqVcra8t99ccAavI
wvXaM68qraB9NJ7txV0gRZzyG0dIvNnvuodeng/OtghKIjjV5ISfIV9tBraAXJTpQyMiL+Pd3XIm
OoA3G4I1E5NW6/Msa/8fIlNZ/FGYRovzrhY3EEwscxMtdjMgvRS/0pRBOPW356F5E9IIN+dOUGSO
wnFN8ZdHCyY0vavfL1wUeH2yj1TaXZ3tWTESQh4vgARXmy6PcGgdYZXbM/QP2+IUJirUZV1QAexA
bPx0q/7v1J0nYI1fYTGsJuJBbZZpua1M0YCi96KKkcc91klUT3IgxpY6BoCH4rzg6q3/uWsxHtgm
K6ib5qoSyJ+oqxz4waSCJ0PhliwUEKWQfku55kH9SLEpYj7bRfjTisgtU6FAVMRqw+mwssYaBqZ3
zti3fIf5PpuqtRiNXOSbF27DEgic8B8dEHlA54y1YowlyJHRUsEov/q1iYBkjlphLjkQ17gr2yWp
8WcJBtJXWnkmpNCbUBTW7pH8GXh+FumCe6xt8h6wVqOUOuxJI0fYiifLl4QiipH/MpntZJXnjNuH
HckgRu0ctBr+spn8MsecEKXdBu9nE1KKyTNDLA4/cgs0aB/GIyGSwA4B9h//ndnV1HLWc2keY83Z
/sQl+1ZATJERgWtcsXpK/vM0xUqDR2yZUdbqCkh+ffXWMXw72Ea3gONNdA77ngNlTPJ1lmWZKhqO
Jxf+II4kZl+NPigp1YIYkiko60EiV9K+Mz3+un/zAjArbRm2TN8KajYey/Cni9SX+TVAbKCCm4L/
AJ2/wQ2cshJkmccsjO8iv2F9puF0S0n18i/qc3MYpvUyNMjlPquWwE7RtwupWUgDdvlfMKBhZLy0
22on68nIb7YcO4fEBoUQMj9NgNjaQK2+LQ3Yw/CgexAlr7bJKPMSvx4O2N3/KAYUJT7jlCqqlrnJ
ma5a8shlEydf/SLzExd2ApocxOx7eneoxi+OzcSXXrUQisVDFSQsJ8jSVPqrb1GE0nZSr0kYNP2C
mHQG9yruURPDYnOiFx/KtFUEL6rtqmtLI+6aKqln6PzBnbMqH3IR2MN6wB09mitq5U6b8bGGjiy3
+fWKETvNaxgL5mc2dI2W1pNI8pUA4jY3Pa7IxnZSVgghUlwJrBdQadtoU1t0DYuUOHblPXqKyVox
EHzeWTC/lpk6ktOhmKLtEck3I3CNcuHnUuMHApfNFhpH3LHpYuEwDeKEhdDkVuo6asqp1Cbh6Ul/
F5mk8RrQ5Q569NeJwob0RsE+93xBcKcS9rzvRCa+orQCKWJjhkvL2HxZtEbA7pRTFUOu4mnpRrcO
rK9UVq2N3ihutU98Pv3xCPtP753GpR75Liq/qTLrGL9efqEWzfqHeB7CPidTDlgOXpm0qq5Lmb0A
YK07+ueA7Gg23mIX9XCdICaeA4riAhIzdPwsP07Q5oQ2MPhT1tU+T4ehYDfotJW4Bu3tfOrahq+u
jgLSSabM0fQ7d95GXjxfId+BTXoKGRmfTdjrnA/Bv4Zl8EbgxQYDNvDcxR8zCI4W+C4oDd2j0N9t
rP7pQcizUpzptJENGepmBMZcd1pzLue4HOZ0XC2Hl5XqG/x7/7h/kw1BVS9xu0PF028BVMmY1U1Y
CFnj1NvPX88GZ1TeAEghZfVTGuW9yRGNt7VL3yFilM0o1Xjqxse3iuU04OM3h6XVYkSzpk0hYaZP
sUIhJ5J+58HDe52SjcBprMhp48P/Y/XYRLsZ/wHZeCU064jKdrBjtSXKRmitBBIxVRXJrKokEHEK
lqOhbbrZhR+w3fcQimG6R5QonbBMEXGRSdDzeNcB1PebB/UIpF0iOMBlT3FkWXK70ojJY2kodGNe
cRYtTrXrA+qphJJgJYawcJ3a23HYdMZ9ASquCp7pd+FghyUsa9dDfewVJSUz6avMWt7Rz8iXP8B0
et7l1V+6K2RB4yK9tXxkp/5Lz3E3uzc48zY3axVx5cexzglgAVdKN3cE8O/Nv/4CbDzsiyNOnz++
JKrQ3lPplRFBHLxMZ52lcH4r1pICo012imeqFob2f4dv0lTD0zsUkxg3/Gl/za+rlaG2DD/MpWks
DdeXmWHRq86coIIeHuNix+QMgy520wUgmfXsUSGPnhw4B3goRlX2IxhBbcZVRpl+xyKmv30mv4q3
1byMATfWILgPKLll4nSYcSkTA9c5rFZQNHj8+g/K7eQa8ghFhwRZCFEKZMpfQ0xEpZSsrWQpz/jO
kxLDC0F4aFp3NQwx+jbL5wMHechjNIb5JZyAXQ78g9EMyfg+ouTmlbbObw5rsq5Crk+G90FmL2n+
l65rpKKB0wYFiWQaeCsb6xlHPf7dUhwqsV4ToGIhhippf2IwHg9VNKsn91egbuiEr7y/oseO4sQL
b2EYkNtHZAeo47mJy15dWNqYNhPBxU88qwObD3j6YR34Pr3owipCgwMWkD7lB8iIjYz/LsNVnXIc
lSBkruhLL/LuT2orJ3CgK8W0G/0PAUIqlnqpyszR8MkoMoc2H43+LNG39tziO2iPXSHk1V5dujBp
2pLjoO/eKW25KNOFUQEc97DT3KkX/mRc0f0oTVibb+HZojjZtQ8KyFb713wNRSYpm8BfGqWTT+26
m/G6vhMQNxoHNlzuW1YLTJ5m7TNmDybiNLb7BU36QoTjR3s5nV0N90YaKvcEDqcu7Vvk84lIIgQl
M6KTaJWg60Z/L7xb8IW8nZOHXlOit6nhV8ixmpOuFN9wlTkO5TiTrxxGNGg1jlHrvnI7sOq53sqr
IRUfCWpWGfQDm1ifGshbHEKQollWnSyqoMjOslxeq5Wb38zxHLhgXkfrKFTKB7fmob9a89hetNXk
bZb8B0kXQ5f8aEoIlnHrdSaIqH1abDi1yznGEXmtxODtRRYBp1n1ekBB6HCdRH5BVQNW+EB2G12G
rwqhqJ6MtI5wJEF12mB3yTl6UhHuo8IoYmhSn+mxf7IoQMOceGQ8OpruC6YA/YQ3owXDPvuQO4g5
RgP2eVTyD1GAgmaNfvE6smm3/Sl845Bgb70hGSflZiIMv8Fdgxhp0gWBO+kaEQxEs3liif4AXrr0
kKmoXxQMkfYK3F5TgcNqlgwvZvBtU4gVFebL8zw305JS7+hZwU6ZBHlXMiTxySTVzM2rILJXsmjy
mC8hj3vyj1OMnHn59cFcdW775aYKhBaadxch8K/5jbX1oPYwRZZDqYeDpP+cWNc2qvO5NBcntSZ1
4gsx96UMG8xi6arj4M82d9CDYeNNzB/We+86Ms3hNUtEFFFXsUafuayDpXtV1HLsQDxoj6IrEesO
36STYsQjoj6H8Q/re5gxseUpNkdN8V8YLHULEbA08nACPoZqp+N2B08rAVzg81Z59pXcdiU/iDbI
brQmIJH41VJd5dx95vYkkYtOD6d6ZwcdUvFuShKe3IZQDkPAwIA1izvLrDG2Y5+z6GYP+r8ZTH2o
U8qBFo/g3hAUWB6V/UnExr1vaMbL1fSV8mXrtrO6y07bX9GZZ/ngA7sU2dLQNKlFY8y3BtFhsQGT
B/Cf7ER+xDDQF5ZUH3+py6lGpOOd3WSQmTLSuQbeF2ma3HjJ08SV0xMGnvjqPVVzAM/WCnCqy+VK
B9bLF9XZhKINlIHGp/Cxp5e1kB6oLX9cKybzgXrqOJqOiCW/hg5NYMj56uC2eVfZTPdsaz/U5ERv
elzRW4iuYX7hz9ZJlvULxX2QoQjdS40euW+gMksH8gdklDPGbR3MRhGHEFSQC+Dp9WuCr9BCRofz
EzG/Xwes7Ylud+5tObga/O+YV5ohsGeqmw0S2iX30iEOY1mpfJtjctBBADgNIjJzUBHzMzPHV75k
BxVbJl2BVr8KI8EkI+cHJruqyOwcHsjOUxwT49FiWnFecFKd+KpOkdLOLcSzaPyxAfAwFEY0YVB5
ju2BjDcEU5e57dNUBp0slbtSaMVNC+kDfxIl5l7OZzZI1GTw4jDmN9oX13GWSkdk/7SaV7FgYtVx
hBfVxgOg1WLXMFymz2jV7lp4vzsGQUDlnbPuKx1qeufap2EvlC9OcbgApzSPgUdBNDjtWZuLyCwB
2RBL9Hdb4pMo2sWDS03ZXzoFWvVb/bilKcs5zVb9qGz0xRqfj2E7zVioAQ0xYZ1COHhvQjOQJ0Df
yDwKJsbh1p6bY/HermyK8bBvq998wR0GiX1kYIP0jd7eLXky5cmMGBbhvY1cZvWNxLzBmFiveP6C
9ih4D0kBz80/pMO/I4WrG3EmPCN8LtrMUG8kmJA0K5UbV3bqjmvBlDBN/i1w3F+knDq7i6wGRbK4
mQb/umAfypIFLgAfjz6PzvsXGbLcX6Jyuy4dZxR3+ytL7Fk7r7hVOhaXv+XZSyxgA7V3n1ZLxp+c
qoEwLI5betylpXcU1me90wf9pK95PAE0a8ReGW0nRq0stQZVAft56iW1jteCu459CGFtpQRLKPEM
yKRGlE6lX7qMnwm/iYQSCsrbMgaMQlCzYmXJkCwHROlLuiB2iJFhThQn+HOO0QOUwKOFm9zYEamK
2O8FCec6brcTLIEMWAaiDq/yngFgdorjiMt5BgxDTkk0Kqbc+I9LrTJmDA3C5987D3sQfJriwzmM
ibtQ8HaG1emMTmH1fdut+lJufQ4n1yO8PBFLYyqxAx46Hi83I4vIt09aNkYaKLJL+Ocu+Nw+zbZC
cLHvZiWi7JoIXN2OyrxOVVu2WB1guBzNRqzvScOQUc/ejWH6nshAYtbwVET9RUnQqNTWtozMRHdz
8NSjWMNtwNH18SuHwuR/6AsDBpZPsVzzFXQfLuM8qdlRPfEbqx6+SXkOOo2f2iqHl2okg9amYAvY
BGeC03FbZiJ9YDwNHfzIUwNZc+6P6uC52gZ9i1iM4aKN4sxzN042ZEObn8Yap7B60qtVCZrUUl7j
kwxrFfhtgWXuntzaGyY7Mdr3pu/usiPdClOdPgu6NxUXgxBWRUgDLcjucfjRvrOC3+INppVw3/qj
6K0qD7v2VhmpsDU+QNDrJuYykWDjoDWArViBU5ASIwCBHrsCKRymx43q1YoPVgtLyytz7mrol4/G
wVuU4bWrg0Ioie72Cc257PcW2hb+5vBkpNDJndfbUi/5uxxb/JEcgVHZLejWXlhu7zpJGjOmCg/n
sGiOWrkOlUeySZtzM6Ql4UtjnYaut8r7ODF1j8lZa8EBBRdugNhkmKP4DAewvrcvxFLEPZ9XIj7Q
XUrUR2XWEC259dGWw1mg+v73YXhtQTGlmj83Xspmksa1RaeFG6WPx4eiBP4dMQJO4bzH9wn3dUeP
NB3HwsdcxtvGW/8JyktMKvEcPptTR5OoiNncFobHO3K12gudZzlwptQQfdcGVWMIzkrE5C0FfopA
/RrJgJkVRAPVFiLek08l8USJtCFHBxJuUsIlAr280wbQwUZW9UbVDTVdiovU+1jmhbwtOsdF7Xp4
8VAL962Lguhr5kKEDrIQiy0Fs3CvgltaVuFodEFYdmz6e89XZuyCKceRG8q7q2tlPKeCfroPxWl0
4shZFzv1QTO3c3qSjtpv2lJQ6pJebHKagfIjbHgIERZ7E7doI5K59gahI3WW2cHQffxfnSxBO4LM
DzPTUcF8busNbTmIX1sXDuJQpuRW9+ylm2/rd1y5P2jkirj3f2x2V3ysi7vAAqoV1ILjeSjgpB97
4ZWJFK/TUr7TD3SoTljsledO1W5Lu91a1y6Kz1c05ZG/Vlg3a/puPrLrc/IuNHGlcVjaxfnZsmuq
f+s4Qv8AHsZGOvHqP67DkGp1+/5+d9NnO5U4G7yRlwTH5RiGKymcuKyDRZVZg8u7YLi7Tu+rXadm
AT8oyj2Ajwf+KQysfThM5cNx0n64B87SfS4lG7F3xEMwKCMFbISrY7I/SNBdPBz+dKc1JCXNC0tS
3ciWaYLvdYtEjU7y+eS3mpDSjZXKwwyO81C8RtRh/v7hG4Fu01oC55umQ7wakfCFVQysLXxws4rW
rYFioDeqVoQWQZP6SgzOx1wlfGbBZ/Kw+6QxMbh6OpFgB/7Swvy/H/vNvMKE0Ta8yHK4uV79l4ek
M3sT6AltNCO4db+chPP8yY4hJgAhvDcqsL9DT4NmialL4ycV8mAhKEJrf3kLzfsdDTcQeoVi2GMs
366Sj3T3H9afSoT1tTlo+fl+rYtpW34uwhdZZC4uvy6w8UwLu5pRaBF3GBsX/7ak7hI7XbpMvzNP
HbLoZVDwnWd95lAegDWXMB5Y7+ajnjrpWJhn8ErREqHymwsfKSwIqC/++UHtHGYFGuekkvvpPz0p
sj2In4lE1CiBIFBbw0chf50xWK8NfGBQo7eCPu9GNPNJxHXB5TGSYIgc3Zd1mJ71z7HPG9k1Qsv/
k3tnNZa9E6hPiYjYXhuKRA1tBSx983rwRFu7RLM1jlB2mDtvsV0OliV9WG3MipfeHQUiDLZWapcl
Ujzo2S+2fPRBuL4GtFDi9XP+aVjD5krXlZ4vu+0yQQtV3aVAJ+oxXrMuHSkUXqrzaoGXhiATn+Py
yFSyjHBXVTBtUpwp1Nzcng2ARmUBnaY8B7UyQYB8qgzUMdagzvd5XFF9yal7zl4L36XNJWZqRw2p
32ukmLTgZMKABfv2aZfajF6KzHq3pXGgpqdT2MQtTuPkElpT9Mgvhj2ZLcDj4w4SWPgP5Ett7+XR
Z/S+kiSipPdDrEws2xvCWg4JUZ7QBDNWBcNQX9ACNtXgGNGf2ELPROxpllZGzy0M69MhHMukrNY/
6E0XVyy+pAFe6B0q6Sj+KTMDwqj+S2AW7c6D3p7XSK3lC12pBq2kKeXrK9libzTzE0Q0Vz4pHNBr
WgN8ZbfshpzcqNmvcZPUA4pypoisAf1KXYamN7ArUmQyhsu9AI8v3/w8ZksUmUA2JWS0fzKfwoys
2sNzca7NdhQoLutKvvgfrTeQLK2wmvTZ99zgABlHAr9HCOlfU7YDeHVt6ZUX9c7KHBJkKU8V8sEp
EoGMYqUZwzYMKf8o8FroWzrnqkkUsoilia4L0MEIpmHIBl97VPTmp01G2XJC7lu3WyPa5DYv6HeA
Fi8FwPj8z7LF8h4wbFV0mNEQfEf5HezzWdv8pcD1exKO/XHdlizD7prJMYGuktgpUTHdGzaWzae9
POtYIkSOSw1m8RI0Z90vc6jrpgGFtqEkFjm1Mqh5g2P7Kzt/Dqw0uOlsjn7GrzEw0dDhSr07FXCP
Ft2AY9nGb9WJW5vws5K2S2jAyCgSfqhkIR2n4fei79NFltgP5pWVGmeAPqU1g/chJf2IXyBf7ngZ
bYPG/M0fEe0PwID7VXdVye+PD/msxpHiBjO5kWxYXZWRw3ASykH/RIVQoL3+pMTnScDcBVEsrNbH
YFBeO2ANdd3I9TySUVWnM44oiq0uVBhdQRozUMTyq6TOUx4Hvd6KVuB/axXtmShn8o+uFihyOxVV
8cBNHJapdAH23ZsuCvfCgdjYhz6gi1YD7O4buZ4ICFbFr0c6H57fPqLhuA2r3iOLEBFdNjBtcLJX
gBAGCqjimcjLm3qf5w25yU2uPJ29C0aOv+r6+p97Nql4MvZILjS8Y0uSu8sW4vi85+f+k799KAaX
JsUvQPtBzC2kYjrUArOt4zO8b51x8uEo4sOzq6d/PelrhrhRRQa5sensxrgFj6pjgLHqa1DLXy4c
+4Z2CuB2OQCF/zFQSjpTvmbY0jPJj/2AeEq0xNjRHoBtxl61YV+pU3d8kuwjc85g+91FBn21jm6H
HEbx8Ihstj5IS9OAcrnEeBLQd4eEHiOem2H1ZHYjatxefoXbvSf9KmcbbnwgJfbXWhKesJoMgdB2
88M0LOsLQQUVPKOknN/MYSyS1AcsGm0Y68coN+O5vsHYZf1otpIKeyLMDOgCvTDjtnbK7+K2U5LP
cZkDGCiM4dHj5KOTdhPagXPpW27yMH1jn5EvjEIPX9AY09OOR2ztbPt/PhaGqFgrUVGDp5DBEBwt
b6TcyFXYnzzPZ6lLyKLRBbGZzrH4VH+PhmPceRsQCzRZx8GurSKD0la0QRlPhNiC+3zRJRmsqKod
rnaz9TJyA7kpjKux+KP7IWbn79aiOQCoG6HnbJFRGRel+qGX0zhnNbjctfUbWZiXTDlqDJ3J5UvE
FVbJdli1IJsN4Jf/NRxWwBKyJyqhYWjhpFrJzNZsJzvhg/n5q+OkmSyfs+XzmVYgJLBR6O1g6a6T
tWDpGAn8FNoYgsARATsYxVFobH89UHZYlMk0/Fo3PR1vNCvCe6DfVi+qylJ8CNU4DLW7cI70+yHt
9DfxKUY7SAAJHAJ51tG9FpD9r0Sw50H5N7IZK7WS2Gnb8haEVhclozwMuUE2tInzDzmyZuKNWjkD
+9GXuuDFd4AW5xsMO3MUFTC0Mfgu9TPC3T/mz2IvP7kAoDe5A32ZhUKHdb03X33SLyAoMFk0rlRX
4AGjW52yUFf7AP8ZjEkKhNbvU9mHRzVR9eQ7e7dGZzhmYdfAYzOwOel0C2GYnqwl6DMe/y/Quc7v
Ri6TtLwH6XrqIl9MtCPUbaxlJK4ltInLgWVC1LqJhQv+7ZKBKPUC5a4hIklH/Nae4PZGwaWgnFng
eO+jCwIqTuE6c0ReE/SfdGLOltb0emMXvifLDTbS8UAaJoiNA9GRf5pC350oSJMEwnDIXEhlQing
yL9GPYyKH4is+wnxmGq1H71kKBKICdu7SaGtbUftrGQAgnOelTjtC3OejiOt7WXv5HnFCj1idy+p
0PL6E4Cnb6tNLEB1Z6TP2bMfassivXp1up3yCMgTQTfMURsa3ub0az+sl8sGqCjk+vCLmuk809kV
BSrd2VR0gtRo9ETqyMsr24cuuk6Qi6plaLPYqiEXsZIMtzgOga8mhR8265Eu3Hd4W9iHfeEPuBpD
j4CGM0o0OnhR4Xi2YRx/BH9ruIqXxgZ65ZG/ZwbZ2Iwa89QH1Cho6eQx0b4Ugi+9HAzhkIBPpCoZ
n8mbRy1gPSf3tIlGy1PTAgQh03v3B31icEowhThDX8qlURTpN+MWvoYMkkRZIo7ecMJmcMioym9a
RDkLKWsIeabI2mVrbBFk8xQ2zHaS1DxtFBjC/ZtigeE5DpttXug7q7p+UNNbylKXEBnR6u1g8HbD
xDACPvPyLygbsvV/uGcrgnv+QNfJWD9mzDvrdIYKSzCySuUw5jnu4xFLjuwOG8HYjmZyGhOA/0fr
FBTNoSMZNsp24h8mpuzWjCblOAjZhznlKk0W+c2LASzzD5TkpKPzks1IVbv/+B+bsKhSLNADyYrj
N6dnujSc0+ztCwIQQzn+GMqmZU7pMB8fEh+peMxWgX/qpQ/4AKkIfuK8QSR8opXGSMKeSCCqU0Xq
Z69CAjdco35I9FIFlQr+yyiym/cyuL16Wp8EdNCObwI6Li++SSbk+LdiV7zglK3NVuxI3v7BedoA
1lLqvjHsfWTZXAF+dlwgJD/c5GIUd35tEIdzh4E2VYlcPrVQIuJ0+oxhmSqbnpUT3p3hAd6gCz4f
NiJ6CuWz8iZoa0bOifp7IUULVgW7YKuWS5T6oL6uyShpUYzNrduxWSTYeCpaXp5SuKP52pYCUjoA
fisiEWoB0ER8FNRycEDijqseTyk9n8bO8b3FIyYIoEyG6qYTDYhEHJNblmfHSVRsY9pKQWkd6vw2
oJPbVOH558PC/Zcz8+2SBCFB5p6lhDt2gCSoUKTKu8yP2axZ8s3/qvrwZ0cRwzrdA5N9DG9MNBHE
dcJSgmGIg+n4zzcHnKbSFfpfWtmM7Aamsefiiw9SLI+HODk7CfLWVEMpRNGmwHEiFX6PqJVlST8w
FeLKoeFLbP6Ie7NfZSQjOqQtCDysKzA9tOL4GbxcSf+1JnjM9CMcgRut6rFB2TCRGzVQNrsR+C9C
pEnB+4OdbQ+j6SiTYQHMRJDoA5kNDr/XoW91cl00zsfsY8khcazPLePZeRRDxF3EZPnqI/R5vh5i
yka5FbNXcxa3r15clrRtJwrqHJCa89mnlKY+n+IhYMnhi9aKcT3ikXfwact0wsMz5JYH6fU3/aHi
JgychXrSETuMdJb0Xbnm3LY7Z9hQdGiOOCH35TEusDNe6LIBP7rM2h0lTH24c0vpCpD2lZpqLr8o
WJ6ocYPs1oq89nEY5nVq2ciZcdWY7tm2rA6mZkYgSBdl2N+44dFaD2mJZjS2en0eUOCe9Y6nVOKg
p572t98gkyynaHRZpCkwQGAmqxzWPzg6c+ErD56jo/nE/G7rW0PU6zV3mwdPLWlDLZDIXRZiK44I
PsUcZIQnUKGxMkWoZfreICcWNoSjgDgqlKAyz1NjRHZE6tgDfvmi6B5UyIeQ3LUyczdk8RcG8TsL
QldBjwuVwPcqFosYLe0VkagQhdWWipA65OCOOmL1UCQl9hwsPX3+7s2iEUZa+tDc/1QeGQz4Vlp7
sJKVxBHwZ8ymFCBqottKvcUbZIaCAyQULRnZ+3WdnTbMB4N+EE7zd+l2wavMJG8X5Om8rfVXjnKK
REGZdC/2AXNdyYt3UTsWSJJV4V5BNfId4BNtJUT+yVlWF+xHH+HOtdQJMyqfH75Q62HYS1Lu0iHY
RHQxGQOQW2x91xc0s8VlLWlTXrFE3izgWcm/GrsnDsJzLxKL9xwZaiqg71fpANa/IOfT2YXzMuIa
9v/Fnzmd+xzKNc2L9IR0BrEpyUdcXDJXYY/RTIPWBwoHXsgTWdkPHhvhLCzPsznmcE0uinN+qK30
uF2ZZbu5pzVjgMRRk+J6iAE91+xu8L4Rt96jvnMwj3FsUQASf48ts6WqnR1tiWDiVB0W5cLM51Zl
NsSJMlRIP5WL19SKnmyWEAhXFxhA6HUQRgt7XiGdQgCg9c9maJA9pwd2KdZWMMQwHa71dE9phswc
bdIHyvQIoFwSuAzOa2/frHKXbTaXvjgv2WLiM3dCeL78zM2bSNJ/shxbzbKRVA0pLNuAvt/CPr0h
0sU1222rvaflPp9O8U1In+tkVnsVR9D1ecPSpB6K53LpCDFSYu/JxFvDvAIpaVstu6tbOLr4+Xhu
/TlqzYQEWJ5YDIFjuNMZz8/M88LvDk/LBi6u7jzNpjFUC2PIFuSiQ8ZZ0cqBQwe8h+2t5NUfgaT8
mD7LdU9/OJHtaw1R80a8NwgHFjiB0TlcUv60BCS4m9SlRgbhV6xhXgYD6opgc8Xs3moGOlZRjI55
auzgild5fe1djR/1ANVz7hQSV0z1LHQrX1Tt/94PuZUL9lraCBTGvaz5dwp7Ra8jRHivMFUeIRvc
IYrYVxE8BrQAUxBxD5QkNUhgyMe5R4ypnMHfnFjIPQ+c4NDv2pjCkWlmGkzlcheyEK5gkBbvMmRE
O5oB8SkG1YV8uRIHtdJnov7jchZyMcIJ4AIKZA4KsZjM4GT/m3RDHNFjNnjdEuZMRaFz+8VJ41V2
4Z5CVqBeMCpyxX28lPWkeGmCxbSTmyzTio6noiUKnjk8b/gr+YYHCtKH1LMrmph6IbENOSjvK5DB
CKBzY6lq4gaChj/CBlH9Iz44GdoqwjA6NtoqIxkSVna1teytGB2ctHLP0fdYrjE/dGRzXGwrEs4W
h0ymiyrlbnOODt+uf96P88M7a0qrDnA+/dmGhWmgRPnBBZwmpUprFz+v4ULeCsAv1Sm0Iyf58+pE
KoiRASjt7W5iYD3IbdNjUQos2bcYQ+dwB9PnurxPy1NxNWweHnyWS2SbR11ucfMUnhxrMJJ6vhwv
pUXDy66nCGJy70SRX2feHR7gqYvGR61BBhMP20j1Mzn//ouJJB/JvATPW1Xa4Lr/q0u3DtTCZiLM
WY9bhtZVbCR7ajwZIhH0/bR7i6VQlWINV42xYloeMr7G0jaDY9x07wuiPQkQxOwLZvE8gd6KGYuU
2/6OdK6IU7EMEW751lD/4qiNT07/QAU6wGWcXiYmLy/Oh26OZuHkl5rpp7OKLzD6J0FpqH7I3iqs
UtdJNZ6tQ/L9WrtR6WXKvehpwyKa05+0quB1t/nvR/VyghkVqloR1EbmhilV95otl7wTXToEXYPH
tLkHh5C54nO4ZaNuEg2d7DhPSICzCj+sWi7lGsfnOMwAV0+AmD5MIJWZiitOZ5mbgGCB+lkVD0UM
AAgnI3W0ntn16ecuHicPVhHgKZZ36w2zzhbCqf7GuWtsvAHWaNLPlEAfGzgeOUyvJIGx8Kde9bPw
3KgLRtXhgLtuwjbiMkfuwDQPnYD8/JirWXeHijv6BL8Lop5fa6+LJM5sDFQ4cuLI8UrMIYgD2rME
Nj2IG2VzsCaisEkHWEUDMsc2vmfbdMh+CDi5342PF79Q4bPLZLCRTS+0k7BKAVv0S2pSSiku1e6x
P4GlWAetBZL+LcDj+ktAL3VSKhfxgeokHU7Q9FJ1h5jz+5tLGvNmo7D7HbuoZQu6LoYDaUePI+Lt
Nt4J/jr67UvSFUDlVPcK2FtXuvyB9g1tIsa+fz0igLr0aUvV+8AP+/E2k6AZQ8hAUKwo9vcFAHMJ
8+9uSdDUiGiBxRiQRiKeeQMkm7zrQoM1Av3OeSLTQjwMBOhwVP6FgZjTSe6mmu26v/d24KaILScL
ULfNH2bTK+HC4bBtgZNjIPFK0h2zzRDmdOufOvSin6d6Op2JCEENtjxwxew1Sa12pToJNivCMLD9
AHb4T1txEpWj5Qs3QzJppVuS2GiAwAuAkREL/otwVOv8TTIGmiJQXUW90pjphOSxnNTUrcKOce1W
EO8LcZ3lOrLK1dwQg5TJ+IYbrzj/ZIZxH/0XBWnBW/Q0Zz0oHNiD+B+H/l5QISkNurD8auAYd/ar
90KBWYh6720WgtFK3vfCfnN6yNqJhpLTa9PqfMsXioz2Txz/8tr6zuQRy0eD84YEyP8qF22C+wjQ
bRFDMwnbBW++MceKT7nDbpwXe8/NHWJG5TvfWweCEzXGvF/CsN6bXvFEclajDLWWi9VK1fv+M0pK
7MUBiBPdwF0JbaX57fcGBnVKDSPjlAunIWiiAuh4H1QyH9MyrFWdS5SQsZEoDLc6UxoMZ/i+6T08
M1BfVXtCRRVZNbG5fzdGcwmqgqbqV9/nxR5M7rapP5Xz4Ht7twO40S5BUW8IST2xE8FZRHySQ1Lw
tLIjkpddQaZB28/2wlNeVJ5ktwzhPW0bvGvRnBf+ArxF6CCja0VB8AWLHrtQ9bIkAfMN5OiVyLgQ
L8ohPbQj1oe+nH/viwJU7jC7vQRheSbfyU7q0gfx2fmDwIQMjoi9KzxKuHEXEwFp8KmhOEyblgOB
B/d7nWVMUxZeHDkpD8NmkHJmpc+NbE7/VEjib5+dPNr/t+b9+DdnCnQtuUHW8/gHz4IzGQNPJkOp
RgGFWJljJgKpmHRk0Wj9qbXIY0Uwfaad2+x/2N48UHVYMm8Xe5ddCJ5GWLXp2RwQ4lugnGZ/vIwy
OitiM6T4s5kqijKQgHYTYMgJHNbOC+AjrliLzXIE+3tB7OSrCZY+u8y6z3QnQhvyjjbsDB/Nak8m
NhRYHvjFYakqmfEgJ5OyCvwcbM2cZoS+wDveyfRH0hFBaSKCofh+Vf9+h9HM3xRx1WGVp+bIjcXb
Es6cqj4Uz62SQN+1hVKFnoQjpkT7aaNZlmbVQKCM/3IcGQTLtOfRrqimbVScfgiBzaVzcWzULCE5
KzqODLxJtxR9JHq17FWoFA5htOLKDvptmL1txL3zYWcaddrcspwyn2aLLW36fHSOu4W9UGk6XjrP
A0V2lMadlERLpT7hzlQgoCMIkKKNp0sVs/zn8ygZ0nXT2AZTlLLXfPZeZXoKHXkaJHrE5UVjOatp
nzw1Tu0uG1t2z3JIAryLmb4mZbrtctnXdg+qghdHp6+1Tk5qaMxA18SHyvOZvOcOujVk7ERvyWKn
SDVleTEdKXXMxO95TAvxcXPF+J4gwN2lW/woMmuGe9DjGoIaIVy7n9Hjes94ELLcACAYF5TqWFoN
QkgTkwW/cdpMts+TGmFVZEVVkJIv4fmE9fhYTlMVdNE9iTncuuLKrsGFrTYL6FUGJfH+qpKasFei
kIysftTynHPWlO2FKXU7IV+pHQKn6q/32rBmtCsVJx8Q3dIE8VVoOTUZU068hIXIBE5GOzeOGxOr
jFLfLOIBw/6U+BtE7ezFxTUn7qGE0Sg6sbmz4BokYiu+d4OkWp2iUqQGTnZn/nHqrSAqNxB4J/Xr
QwJQ6oMhCfXHpJplZjkQMF2ksbLYA4eeNJ0OYdyzDt/Wh9RhbbVXbKEO9VswGHkakiurJwqAoQqG
nsx3qUa7v9ZDb7FCRQtyDGfLoHoK3MlcDDTh7WY7AT6sj4Xl/tji6kPN6fI0oW6UyQ5NfYY6UTWs
db+Gawm7hJyl92wbLqZSa8IcCpub685vPpowk/dutTP+lDaxdSAG9FARNA1e+QHB1nhGxUCNBcR5
94T7ggXz2SKafJaqC2Qc+k+tOQdvMf470VVJjusPvpf+jitgEuBEjZwsShZVeEtK3PLFYXY/WLXI
ULJChTjO5SCZxJSmQMSOVl84cBZSOzetY9U5Svtzkf6DNCDz8U76KKd4kHSAvZu29i1zYRST+qx0
kPkVBQMk7n/1EXnz4+2JiWx0UMPFJoOhTpjA1l40eftpLDy5zqDvcJZ9IAV5L3E/1p6RJe1WOm/J
jyeOq49UIYnnYyi7Fu4X+qpq3IAoT4FCnip/Y76r49T44i7NC0euOfVYUNCceMpmxMSUa9/8P369
egnjU1nhNu2IyVo445Gfap3PYHgDkmotTgEr0dqr6V4UW91oxT1lENT9e8AcZvO6shsvp0Px3ogd
sBnwnOY2h1KpaCK6HK8f6mbvyiKR1WPR0ULzeg8EVs+0Bg1X3mD8GA3CAgt1LPSqQwSp9JJMAr/6
JA1fjU0UKDHDi0lDarO990dADlcBSdSdb1Vz2+vId9Z57PY5gjc0HeTvyPYRXpqlJRxt6u6zXmKF
fQW/6PZDpus/kevS8ckwX4uaq5GZSZxNaTQ2WlGVttGtCoVC2PjYQIIocYAXaClqt67mBPW7pO/u
yT61bJemDciOeG2T2U25+eBvOsv9/fFLpQMUDGAkldIQ+jmuYvUrE6ScRA1mEbhkxI815kFvomzu
DseJnrW917/zQjhp/nxls1QdZQQp9+KhsLzKprODgPCKheoD4wWKRP1xdwRC3NR8wF2iWC5s6jKv
GDOZqXlRdHFR23tEeb61sBqREK389QhvYWHn8bObntmXUJoBLX63Z+Ky+/iBHttc7o4NeOq+5A7r
KT7BohyVtoxZhgJv0Q6zxO1m8z5aiwYO52P2XSJLq3Ffs28yeFxFN+yTF321Sm3N+LoxLAszGplc
6kd6riQHeDV6kBT1Q3vyN9v3YJg5xIU42gq2FQbAfhEtQGhvAo2YmdBeY+yecLX3KsNe+8iTCkLz
HcK6/DutR6nYEU3hBb06LvZbAxxWZtdJZfzUDg45CDIi+UntWujget200p818IEK4i+bb7kiI59K
aX4eEi0a/fXJRPyn2KPyIFevv71P6M6oYRIP/c2yTYsDyhDHB+NBGFrVXuK1TFBTvtTRZf4i0Mlf
eok/9T4yzsRHTN83D2YAqUM0hoRtZArdegUKSdCEVjeKAhOy0YC3ccShYUjm4hebknaGukqoZlE7
nxyeLwwqKxnQ6VrahbWmXL7bSfQRpkf2I2a8NLESX1ED5P7LvA50m5+/HGecD9b9/E7NyvZJbWEy
FgNePHe1dmqxciHOS1kBrx7ocZ56JPikxLVqjRWuefrWmBYzTAdBQM3+tfwUH5pah/WmaqmzICWP
9eXumOq0Lj+9h2tvLK93EsnMM10ZZMErdXuGBpIEzQ43oTE5oGzH5KonQShpwxNLCja6mLvLnXZN
ddPs67pAMKbqDoYmVazjAFGUi9R6Dz2ccCgDMgCnSsfZm+ShZWG2+eU5kOCmaFCswu03lbXLBF3j
VoDxgaUCUxB2ol89qF8vVoYvCq6lYpWKrScBaf1dX8YfH2bAeqhq+SC7WGPyRxVYaLZoiu4Q6M6+
YQviOXrG8f0iP83YJQ9i+3HIQAOybR42jhrQ4Xvs/uQjE8jGh26eWEojbNG9j2bqEo6aO9IITcMA
T8Jt0U14wDjPnO01j0LauZgZpXxxHiw3ArUuBuFdNEt6uXb3fZAn9qebiNfzNVMBbZToGCWywzB2
uBf2WNuKIZncFb3XzuiEerIi8xm1OMYPbONgwHsqqNH+C4gXAO7yKulW9g4tgGL70qZ4wJ1ycQdl
9SBUkyIoexhzERawqSJ6RlG0FexOpzqLI2gqkds8VKfNCijce8UoloY3XbTa3iwd/g1P6CFxpRXX
mFMPFInzIo9xFkq5+YRVCGJpmH3MberZ5FDf3iJhkhvXYar+vTc391zPGMvyKkwnV37iehmIKqRK
jauc2kf0P1jhIbaZR6ZdPdKNEftboavcwSLw7drtsKfcH1OFrJGjxvnAvbk6EUDpPQ33UCcD0YA3
ZHpTpA+d1oBKX4hemxRBgT9RSTfMCAplaLLdQrptjtKhVozjn86wwW8GdhSL4AIyypwsGy8ogMPB
GsiFgEb/PNWmcalC+8TGsOFPX/Dzb8uXirYlGNA3CfZSNPKXZpIAXIERDi+q628X+IbwH1ijRMF/
0kF00xB0uC2BvGqjwSZIm6CyJ6GDnH1NQBtWGZavGxWuV+R3C9v97k9Dx4+vF8esLQFAD4Gypp7I
g34wgPXiY6HcUJi6t1prBvKNDJoIh7o9B1NW6drTmDXSL6sInta/8+RDc8vO8lO8V5Npi7z9/rTF
5ocW9bqEkbEwT0kkkX1smhSeYEjr9sy3eGNYLeem/z6u9P06krurF89pd5s1LMqJT6tKUunONWyu
/z7zcIypciDoKj4w30B7AypO4LosZ1UrGsMop34eFD95eSrzEbqXvyd84JhR5QE40VpRUy+IJ7AL
rBZK2dxVBolxZqUgMZcuQcOiznSkcAcBA3cjqQkIrVswyD7HfuvUh7vC4eKzKuR6H3W9ErI+72yp
AlK9Nq3+Z0Soq5q7VjNfH8APDTq/ADnJXp1Qv80MJqcIDAUvP1YqrQU4Ql9rJzQ7/4NczGqVPwnd
hDy9Dx6K68yHaK3hoYhjDsEVY8zXcyl8B9RQA15padih69qXuWHsPEs6OQPCR7mMuDpkqNBnajR3
1SYAldxqy2HmNUmt441Fe6wr8akn95J3L+QHjTqGBwQhI7q1MFjH46azKoB3sbTrHXAJfAuP6hiJ
AaMug/0Lkrk4xoRA0vVWxj9sYC1xdho+M96J2NfSro0Z55qSDDvn793sV9A4Jflh/kg4bAbKRwuF
jSl0WYnyl2enisgu0D3jg3DTpo/bfHKQNheuYatKZDBcgt9tcZn4s17t32pWhNoCbgNGLb++lPWM
sbw8TJreLrWpGBAdWX1gt/sqONZs9sYeNZeN5BkGxChnyW/GM9yNrAZOuAMGRv9dvJujJsIc1O/k
76W1CLRj8lef+6EqdeOdhnM7kCHiq3XEsrXMeb7rGWJMXjRmyc2fCLUy0mUqhRnnUd+osWDB5J17
LxKeYrIbCHFjs8WALB5EFn4Zkiz7sdI1JHaMw1wIxi4l3OLCi4cbxgXu+54XowEH8nf+mgJHxw0d
xkXzPnUU2+9fBmQNbwJcY9fUH1iqnZqVWwC1bflza4/aLiGI45XHhFCljNqJ+J9e0AsKrMF9sGH6
x0sCB/pzX3W9q1uImsAxy8uwLMMd75HaSqG910CvbvowedwAfV3dRoK26wBVf4GoI1hXuAVCd0Je
2OaOmSjaIdlc4WctN4BBo5NR9i4b9vTABD7y0pM5pgKVfGklQJnAUsMHAeYnDkTrDVJ1MQvXM/W8
Z/KjRh59trbsovjYzakgi/udnnft1/1ZCZa/aC6rLK0tLaqbtFy38MdNyzzLAFwOYh9wveejes6A
14CJc97lR+95zPa+dtu4R0tW08ceKF6n9NKur3p/zIdV43rRis4Q9ggw4LWFLqmrVgTjBDN+1OL3
/cG+qJdWVXn3dKQnivquaTmXixiGC+gqAYVDVkOGrr9/dvmic65RDINFfRe74wE3Qeoidd10G5TA
S8ueBFB700axTjrASBXYpolLj/LKAEJfuWgDDASndELt1hDReHvyKvbG+vFqByM+TtIlep8OvuUD
s5GX05zDMF+o6CqsrRHubLZpxgtswTczStv5F7u9zZQm9ESx2l2iPLnr3RQN1gYCsLmg3exvrNIx
1t+Zk7E9/JEQSQ+AdGOFTEJCx0EVqg61RDhMOJw6EJglOS/blMzIHbYnNJuQ9F2HmI4I/QQqW8p+
oq4H7rEK2w9dZ0Azju3LZ5SsrowKbfs6pVEWSPsZFnRLxC+0lm1jNnwofeFnqPGsPto+i1yd+0D1
BRYnH0KOAWmvHWJ9aM/DeKZb9RRuSlVWaBWjFiV9WLLIbqUG88qRH58Nfx0tlPWweSMD52QQX6S0
C9V0vH42+HMAXid0nqW6nOocxnIctl7y7hMMXkbDvsbXTYV6aApUtdvSjyidPTJ1y0MVaZDWwjoS
mlbiiqvl0VRXffOn4W+6X6MW41Dc/KGCfHETj9vpVREM3ZqCoab9R0KcyBUEliUt/lBXeEOvrGta
XtsobPQMAkSUbLAekwgtko6csDJ3g/pBvtDd3mzS95mnnoIGg2zLsWaqnKR1vFZ/n1q3RnWPdDLX
k8auZ0zZuyS9ojjthbXNvJ0kGKO1BR8ycWxApKk8TKGt/p5R4mA7SEAxHdFTsPVu3wdQyQtNTW7K
RwIpXyTcPSIvyPAdyKpCEFkIXsSd7PMFiix3mE2uYtsJ1K+LKO6OuRoa6ayPnMdEBa5DormgYVxM
Ms8caUBTy15vwd+Fl1gxzeGZm4DyIp8wb8udqeBRUdpmTSFh/VrUXs5zddnhSZogJY8XuHFXi+TD
3mrt10V6g0zvlu5e9+A7DJftFk+gIo49aY8gdvO9cTe0Nw1k8UNgghdlsPGVUEURQ1w2oloIo4s8
1GU+F/bS4bnGEw51745k6JmttoONxxsjhCVrOTrNFbyXCodswmX+weglIfC9px2RTN9N6ubjU+Au
v3gCKqfEri5YjNavFJvYJ7MkT77yPF3vFuO/ZSKmEvScky0K4azIRTDAhoGgoSxkYrchzJqpy6zU
Or7JjOWurSLot2+miqH9eVkKdyRNvVgt5RUm+vjByrQ8OdrnkhZdsxa/5KAB6aUHzPhlEOGQX3HT
0VGTQTrFxaXiBSZtM2O3TnnuZY4BwoNBi85tSceMgf87nLu4lsaOXl6v2YToMPKHOVbnVtGjHBMJ
4cINspRLt5KvD5mwJ+414x4TCDSdlz553AJ913hGg9xl5ATFdTGRj6AUVVoURyTwbz66LYcStH+5
xGSzUWhHDL7DMQ6TYz5Iwq0DYtadPd/kd1K0HrDc7GOr7VkTbHqCdJyDNznIaIfRVGpqu+2WtB0R
E1HBb74T7sx4RBf3GXvVq3xiBFztpowcN0TjcGBkrOcdyEULva7KfecxPW18YI8mpnfIyw/ye8q0
SlCrO1UOLkjYyz1N4li0MqOHDv+rPDLPlphK6TXQyj1QFf8o/9PWO+RZ/ItJe/k5LUPSlvYsnD46
rUKxE2L49PRGx7p1dHrtTR4Pq6eubPH4UWKJUAmfFbSjyj+Ow6MdPY8G2Trf4oI03PsYd7y+SCCy
PFgvUnYTGz82XVgcywClTGlv6dEnQoAfU1DLY1YnRZ/zKFiy99548+gLhD6wWMAslu1l+GvGvTB5
XheOHMzVovpk2UGK5MmE+Huw6vvjRf+uED+fEPM7VG0HwHzzpkArN3mf20IYak3FuLmeDDifa2i6
HcPRiln2wvglyvfZcsp5bWs4xYi6asg9THDDt/4ymjcLd7+oYs4IwvIgyvmt8/1RSaemTI2ofLI9
iuMhKnn6VxCYfyTacxhyNxHrTGPopm7O1XtfvGO12Qnb6TQmWFa0XFwloi/MG0L2Wpk0LdFOjH78
iTXdxY6VXmAc6g80ZZlk1nnUNbd1H9HKFiX/J5b1EDlt/q+4mhPq2JsPiOSZ8p/AghXSulLhADbc
UJoDHoE4Rvc1hrSJNbIeWZclCaPNA05w/ebKyAbfn8pBVT9guNuowy+AYn6jIxZ4VMiZb+zJt99v
ikzbf9i93IPvY/0/SjWszQ2uNbLZILk4eMsab3+mH+IQQkEV6fmxa+FQ0Z7BxsPEvC6f3UGeFn5X
D3SPxbee0lzfbRxBPx6zNEtYSBHX1CMSUB8ACAM9vPhljK9bnBslyveto+DWMR2vR0OxWBuRh/ro
tXIu0PhVDF90JMBZfpSQNkBu9xmiwhXGSqek3Gq37p+bpFSMrjXSS03LfF2BHfRksWVj7Cijf5A6
zc4QJOVwUUxoblo3KbyPu+FJiFQJMC7jFMpQedbDie2bwGKpW+fvWTM63J2K+S0KbOYOg0XHck+3
qDnfAHVloyY2/fEs+PfW5EQNNsHNP67OaGaDF6cega7VRtZQs74/FPzEXmenqaod2oAM40Nl2uHV
rBLY6KuocVdWhP5Mfv+UMrHlIkrCPgnJdaLQHduSTpIM0BHJDhwzdhUiTmJVo+HfdD/8CE9GnA7h
CfgNLF8X2xvR55j+z9d8q3YD7tybddNbpTW2A/f8RY/9cQO+nzrREJzT6be8Gt0bQ1FZoH9xlRz0
qi8GA9QG26LGbLMaJ40JNKITmuDLmYD98fiFDRcIcazxX56wT2ls9KeV47tk4XtzC2b+13dlzBA+
5uJxJyAHnJrMhfrjDz6DoqIBy7T+SXgDu5wa1cGe9hX4X6mvdSUH/X4/cUzbPQEmL4PGIGmelZan
7ZMSGHdn9Aa/xRmpRcmOp6iWl05fF+zt8T3yDrpoJe1N/zG+AgdIPzR6AeA/RvoYK65XCBXMXsLl
b6gOdYB/mNbUdQhvPAHbh7FnP5+UHXASboZAyWeLUBILYtBL9PMi2FXUbT7S/9S1ZB6HAWgzvTjk
EAxf66S9FNvMoguoPBHvqo/Mt5YTzEaVxprOYqPUp/55zl5hlPpQCS/yYtCm8r3N7IOAa/XQY3y1
WftGeHSafIcWJYNm6UJ7o8UNaqitvz00w7iI9Kinic8ZFibdhB9xNj7ZR8qDuQNHvBYKFeAAVPo2
Y8EpwElFm1Lj+fc61snzMKrSY0AM+UlsgPBgS87agRckIn7lJyn9IAYZp2rvzhGpBJPrNlt7PzzE
XpW2X4n4+wf+TvoW66yF63BdyT9ljVG2pkCZynpV3Y6tiLYAta9MZhpHxC7X7liHPhB9EowmnZ37
KEUiQiiLm/gz/BhMNkFPAvvLquJ1bHmiBF1VTJlWgehMjUxmHveLu7CK6r0eF9gTg59Iom1FtFiQ
fCIqE6hssDpSDYaql8dRIAwX5Nv58xa8agnbM1L/V3BbDA13pDyRSt7cppctSpcTapF/Q9lfl9Sc
iKFij5BMuIqsgQ1wXwVrD4ntkfqsyR34OK9unoLyCsqx8bweiwcgDDjOtEO1du27ER69FVBu7Oc0
5QQJBGew1964nQtTkuyALhmsgv2wh/M8U4NWLaPzZGVtvwGBVFS52hPaA+ZpaD/JhHtBK/OXZwus
8Gh6pZGP5DQZfJSi8Ye5i/N15hMAnahFNgoO56yVzSL4piv9cOjn8KbUzAlC2/vNQF0YNakiT/rG
p3xJTh42CtNsjXfXdzbycFaiuCKQdSRxH9XCXiYwXjpcBKzNcGbOTv5/bwxs7mIqVz4U5/P2zvUv
R+I9d12ddDr2ICoc9fKayz6Pmisg2Ofl+sRIy4Puq/AoCACJT320t7KHcFpysl+5tuQhLv2wr/Vt
M1sGpHtOmyNfuA+jZdymyvxG10FtOgm6sMWPZQctx5801aG9+27ch9W2CeoZH7RxNVuYDSer3FOB
D8uJIycM1ks91Gqk54o+t8K9iRquiFbf1dfa/PTtJDMyQF7V+5/8lr9ur+YBrLvcILubMi9y2GTk
FGZvTcfKfXcqSJ1QamkJ50pbXiAdT1npLUZRgx4JQo5yApnttQ0BhwfeqZpkXIFdBtkcPalCNnEw
BIhrvyGov52keiOh0k1DuB3dSNMA12P2Kx3MT7dref4pc3DzGQUJ5loryLZfK0CzhIlKeJYZJw+M
Cr2+FN3Qv/kjAT4apAdfQWuLEMYLh6f4Rpyo2I4QVY/FmIR1Qd9cgJyNz751xOaTiNxvxLR2QUfA
OYTwM9fBV6v86cwZTiG2NuHU5zJLuBH1NAXb85TA68V7bbwXEOeiddmHQzyAZmVRYsKL2hE7wo9f
lcQJH3FiZ/BRjg6Tkw61CAxoC6/JHUfZXiuIFcpy035YQ4CecAxGkGauwaY5mhbsPEqW2HS4x7cs
rBMkTM9XUak4r6+fjzknb7ITAgu6bhmvM38niI7dJv7bjDjWFb7yY1Q/tbsnc1WdYisFhWWlfJJB
ou0ZgMEZv1umKYGiJ4i6zKIOlE1fqRdHNlM/lGttFrKdbmd2hGSA3HIjNsOM2QjYEL/MboFFx9DL
9O9sC8eE6BRDUnXj1asshFRyU+aXmP/V5Mel8G3+tfbiTJV1roGRzBTcIJNzPr0NHu66bscm1HKR
NXVZfsBneJw6oJz7iqtk27e07nIqA/3LTO5slJ68/7o0AQFzA8VGnSs1zcB7AS5C+EEx13hWUCIU
LgKLmRdOYrXpZhIy3LvEJRQp+vQyc2jSJoFoEAMNxZEALYDmBmoYFofk/x9fsppfdSBBlRwITwru
DSpoqLsnZT1fVmIzMU3723VfTSyDRHgo+PKh6rnQCD0KbbZoAHwmyQYHUuoIzNHk/Ub6PdbPFtRe
4gCZQa09uUA/wZifrH6gYqyuJ+UwPkOwF8rPCqcivUb9aSUd/HK+i1yEiy3Z07KMd3P6z3Bxwpcf
15C22Y4gLA4MbrnuS2zlh24ebYO0ohMVcpEAJXEu22GawAFTo3hSKYmmVVXem6vFwWx9s3P/SNm0
PAforhC8ElcnDn91pTzz97Ht9lwy5A/1lXgQn8pdxgViJOPsOIMuPERtoqqZQZPC6vAHJ5gX2Hhe
JXuRGemhzhmRTe4KP81eaF3+me2VFBvyTZZwYGoUXu2184BmzbKdLsTFSlyGrk5dkJVRM4GAYFDu
2UEMnSX1bwH1UBp7u+wviyqR1LKetSfGdCsYKU0xv2YzGfEKrLluYyL5VURNjcRjmNZupdCqTNC0
mMcgevuVy2XyToXOhj5AmtnfsAYcTLb1V5LCHAUtif3rJ45rnQK+JdHPHqw2q4GHn0ePL95mzMk7
u8h9rgGb8L1oO+27Ax7GoraBM2V5mUFsGOExFbtzQs/49fRLkuoMNIxIQ2QMesTvJbLVG6YL2ZLa
ZvjMKuVEbWrutfrLkS5aWcxiSDknRMosHPgN2tacmTp5IwGLN+iAQK5/+aYDFujpn8bZra8R/+x0
HgSs7h6n5AL7bzW51VgYNzW+BOIgAXEObp1tbwqLwlu/dJHCc0bGDRFA6BQzc7DrUfYihK24jOUk
nN2Z6w0HJChatzLA5KKpgLYg4+Rga5BMzjdza1BGGzfR3s7RclDR8f6MFF1hn+I+HdgoJo2tavEO
sUm1mCyoyHODlGpGOD+2zwW20RW6vGyX8CDWZfQhzv84MADgSsias2+MJ0b8m6f2whIIDMeZBu7D
7LMeXj60RgWxGLkq86lBFPpNMaa7nH1pZu3taZ9ckaRpBIPGQcukqAxVVoZBKL+ebkI2VBV9Tcgq
0t0O8WCeK1kT6V8rUQZc+IByIKBr+FhMORiW5wZYT9mkkcK7sXkbAHJiVbxNPPSp7dBTnH7bWtJR
b2/KETlQ6rKPV920S7VRdSitRL9FleCIfP4GAMPhtM3GEArPSfh0kuNUuEf5vTfHccFChJyo5Z9j
1164Qau5QVvlBIbw+jYjViyG8ftm1qd35qupItmpDoO94EOUS9J1frzFzTOCS1PzXG2Y7AgcNC2O
d6iF0ob4OHSAfF2mkkpdO/kXPo3IcYHvn20Y7q8R3BdaHQqexUUs7CJn9cC/ISR0PhyvZuNlDY/O
K+c0KkvQv7VJTocHEH2fKPWZr8PbP/2hnVcjuW42ToI45zONbozkn8uXzmHXh4X+Y1iqxqTYHx76
xOY38jJvRP5B2z03F+LLuuaPjuaEkZOFV3FpvGj4janORmhBqwNe7F6TVw0sCpXz4dJAmmK5EZcX
JcM5sZW5iSJJsOTfLlGr67HKlTQeBS651RCi9R9wUTX3nMK2k6dWzv6Ic8A+MIIMd5R2ZLu2EJ5i
PdmrU+hJFfwLPfxNLZ8ue0aTpV9IvIkAaxNCb2yXWo65TFA6Y4uq/xAH1BU1S6dHst7AXijwoOXM
smLuPrfym6kwbAlCpZj8TPxJFl8DKo2+B5qW9FY7Ov3LFZde+WgQfjzSGFkHd4/DQrOdPAbCkEJq
ycE0xBFfQgWc1fGGDCAlG85S8xSf6YRZ7dQbDyTCc3cDc+DGkgUB5Ra27PWiPxqJg/UERgASh3kf
2iEuwYQJ7W7YodZBlE+d8I+kdiFs1eccElwfKclu79PKio6zdCuKCuUXjZU/5K1JHeY0nyWc7sB3
Sn/dL0S10f6NWBydIJizD/9lvTiRiDl+S4TQwyDpskW4b6gE3NalY91IQfCQ+fPYXzjM9BYk0HxB
kuQO2tiJJ9w+WhHXAVLJiLuqxGqdKEf0y5pnVbE16IIkhTR+vhh/t0m6gJahcFwoT+fgcc1lOD5o
pM2Kt7oDlcTF84DSYWzpxG8tK+bBDVvaq9cEKM4IdegqguCwgwyDufm6/tfYVXkg3toyLsl3d+Rw
uNxTd/6tL5LIzaotmvjAKZZK1zASoEJre137R7FST4z0cCMU8CtcT2zGdVQ6FzxWkRYY3dCOcTuz
rdUWBDbILL8+IaKUCAokP2emXiXdaWJcC/7yki91vDTaOn2dGO7VTWvV85VEd5B27hprCOuVRs/9
VtLV3tWToh07AgIS+Gk2eUAyDB5Wk3zUwBzh43JmtItQ0mXfx3q2UlXLsFdiltsnUOUsThA4ajS9
0nKxeogRmDt2uWsxKV9ljJejQoHHe7R2nOqu9TaD6bux/3IAGXQNBw9Iwa9tRTVK04DfJAyWJLIy
qaNxLZiwfbEOZ8f91TcaKAfqZkEeYepvKcFGFkIW3TTfNMa2Y0Jlg2Lii5UFBm/VIXUBvSE6ccZK
npcNwmglNd3GT3mNZPS6i4jgnT3bqRTimffa65AOfE9FDqN6kKMQeSjxW3Z2QGt16HmO7wsOxoUb
jyYgpuUEWo5HGbFvRmNnQdCEfOaPq+dEwbeD3AewvmZNnunC/hQuGL0204P8WsVhyxAvyrP6OQ8D
4iIpe7+JDwuZybK5d41wBHYKpCn44Jv7szip20THJ3vEaTyS0o8iaNqa0qWI+FY+Hpw4SszdkCJW
LVP12zh8bA8X9rcI6xPk8FU3W7+OXQVCJAneMlfsOQpUS2mQcvMptKxqi9PGGAw/JZh4bzlw0Pyb
scFaVOZBDGfNBe3t7qpOdqVlmYg7fii9pxxTGLDphrfr7vCGveKzMjVF6u6ylWRwdb6rzDn2Ua7z
9q3+v52VKl8HHnPJcZwvbms+NYQwdoS9Ya/KMaqDXh3MBhn7+XvdcyTcP9pNrJzE/wJpb//ZvEju
zBI2vF0kg6QhGGTsRFw5SZhFuQ7v6vx0wbH2IciQ+Dmqh6AVWZx0laXf3N/921zjbTkHmUERM+LY
5GpyRPO9zhwhdY8dWyn9rzaGOpvvcA3LXCrUlshOVO6bvQMd/OMOqqzpJpoYZEnXM3PVDsttXlGB
Nj+J0Pp3kPHvKi/Z4BZFt/yEUlWk0mAAhbBbWVQaOwvV6DryBRtJvh19b71XkypodTJaTHdURsDi
lxT4tU8HpNzoJbBPfLE4dUiYNu1QFSRpomlhxQQSMc9pFaiFyoaJ/8b8jVsaOKsSDQIWXUciLzPK
xCHhoJabc60Cb4BpG/AsETYzcmbCgm0GL6Ib2RVlFLYrrCH+yTSCAT8hzEmWOSSZH990GGtgHM+c
SnWgNsoxGpJaZOlSG800A/bA1WvClRNSmQeyP6liIgetVOttXUSSQsW2sTl4WxB73Av9BrBtR6O3
1/iniXy34BmLxUX8n+4dwskcLTjoLK2hWitfodZznqWnsunDhlEKnzp9ZvmMPIANa28891he5wua
sdRdkmTo2FyhveuEo0vrdfKeuA69lAJugjeD8fgiDxZAwxdWcLR6eXf6raCoH3ynAemJzUtGqEZK
TuysBpQmMo0ioy8YhquWNLyojsBHDxFNqGREjgFyptOwSZclvCydizbMfLpTXQMf1OzOYlf5ABoF
kqv5kTuKvAiADCsDPf20DKRlKg+Od2Zpg23dRgBCWZjCk/8RXcrFQqg9QjmZHVWF9zS7P3JR0VzK
2MvAj0lFL4DoIopgJcqQizcWIVsKDIKwAWo9nJb1zxwkkhSz6tt+brW154MQ4u1kbLnr8iU2MiA0
XhW/E7T+Fdh1WTelzN7PymsMngte4fAGx3qSNUsAPXIc56d3zQQqT4s9w3NjurYg9dpL9m+z2aqj
ruOacbQF6hx3z7WHWSy8/fet+ilEnPwjZQDKDVgC98aOkr9HaFA2oh1lRfaHqb0siQLoC6wuWYTN
40ftySvmkEFa0iFu8cFacPwLOSHwur+rMrPKEvL4xu4C05pdAc4ymtvZyDTHsfQRiDBD6jGecf6D
i8MUbamU50zOgWymJssF/ekv+7Xk2b7ZZ9nOY+UA0GL7ZE9B2b9Nb2gUnYh3X65wmvfcF01rB3J6
EZ58LkH04RgBgGWOJd05gp2k47nxhN5UDJfXlmiIM62OBgCd6qlaojOUq7410yJk/lPlT8z+hV/P
liJydDWAL+ucUiCXguxkLmi+upOk0fLskEeSzFygZHnLiWqLC6Heu6JFhxgIrhFk0NZB6bxni1la
xBw0W2cVi9QOgeMU1b/jlwBt3ZnjQdGEv0XFrnceah5LMq9fp6sTAR9S5b8CRKUQ45pjl4dwKVvQ
Q+tMjO3L5cnX+HJcSwOmsV74H7j5HxBJiKGE5oqyPEBO7Qa4GX+ShRVwnGiWmrfEH/pv+dOxOZQ4
6DZdHai+SuSyyWeX1PWu08lR5dZTxnOQEr++iEngGU0oOD8bF6heVhRZ/I/oasONNFk21f11AUis
jjBvFX7DR2NkKZyZk2qG2vuNplhKJACOqNbJLUF3TTkPlc+fDWhwMa6snQ1n5/gl3QvsugFMCM8A
8vxu+vqBniSMaurmIDiUtkfM3V3kMdYnaWqzL/9Vw7hBmBtpd1qQYb62gN7UVMVHFNW+/NY7XarD
x6Lpk33QTHFUPume0PQdY4ZAH6InkdhP8JyIV8Hv8/5hvi4uyAPu3lQJLCaacXyK04TDfq8Mva9j
OaA1oLbG8/6lJ7YQtE/aWAioesLysuQYeG1t1VCP5mMZJlnw32dieww55nt8F/QpWNOXSC2Qk/IX
W/W769OWZnnavA7cXKNcqLINFkxYtouinYtoNwch3ZJc6fvKlyOOjPRcQo+VYlIo7O3JJmpD8IEA
ceaB0623eXQory20ei7fbzXbIG99Ar2n/4WT+GNO/VBlOzoKG/7hyzZW76axnN+C/HEqmVhF01GA
DYhobIOZSrkGoUoowAwMh3PQNLmwIl3pnUrUNtASxLsDU1W9UXNLJlDSHh7UyF1xnTMWwU+12Sbe
tKLW0TOKWNZSPFLLQMTOm4Y3WHqkb/IU6dFRw3DwLRv8Ejtc7md7QLALvMwEkmaJqiTL2X9m1t9c
RLmHNEWlTfm8D14SsojfGMZ0SGx7dLCv2BksMVlFdXQYdm3m+jHC+BDg62BJNJSajK5lY4qOKoDz
NlXqYUOkJ7uXRBW1x0KdpgJnY1MXQwRCzNnZY4vd1sdb4v4oR63w2IuMMQ62wuCdIXwmY39W/Dk+
ID8vrs3CZaaYtziMAnf/5+yzJ0ay9zNHsFy1yvXhR5B1s+IjM/Etgex1eK6Fkvrv6h96YAKeTvHO
ZNNv9vz3S+P9q1fZOk1oHvrph/eF7CZzShlOy8PiLY35SQ1J7eOlGZygW5sr5RL3TAO1OvPbA3sD
LqX1zU/MewbVHIgJfshNAlNRvUd0BmYf+kTEiMEl589zLpwv7xkEMVCYOEAhjM8qd7rq8m1uPIVD
W157Gv3wY1Ym9Sd5aQ5bTkm1pFCON2zR/6I+teXGI79QbLdvlJQhfopzelv0r+vzXjvPCylxdPnx
EbuZhqBuC7cHSHvILXIy3zycfKB/mylJ5Hy/mL+Eeuikx5H4TPnns1RuOKucHP8ySjRmACaP7Txx
DlZK3ohtWCpCnjaws4EFxJoX0+B0v799XrZgCqMHqBkIInSwjrnfbe+5DEg4fRE+fcn0GRfNNwK1
TEbJbMpUthFsIj13I4HardokGmC4SFrXQssJrBK7vfDYclfJlDERF+nPWzHnDJyCY58XSE6Ti4VQ
PboGJv4jhf1A6anyXCxHMzLMImxuRiZ/RKEH8VtJ8gQPqJhAYfx8U79JkDaeZT/Fx/nFEbFle83a
16AX2H3JVO9qwCyNRLxJagUvyhgRhWN3MYMo3MZ1FIkygyNZRaarXsJIEf002uq9M60pBtQA3s99
jqRkz38I1wGXGCOAFZq1xiW02y9Xxs26VRSWJJFYSoiupCEH/F7oxwCLT8dWC6THZ6SwXtwT+0vK
MgZilAcLgmiivqG8XOVwhBXF9Z5To/PEGXzbpjVN3hcvdmm6d+f64PEbf4cZRALJLACIjQFZp9m7
yURUBpWHHJyxZIKw3eI/6jhGM9pOySeu24Myplg3A4XPfHchWIjSim/ESEud+Y5TA9PfzD9Z6Qtk
7/PdDCnga1XV5wBTCQmbfbo0WEkQVxzc5/iMlejrHOxttW6Wb7tf0wQgqoukotRMKGiK0REiu+ub
FdjTggowyquJAkscKSpOF7qpeLqOiA47enr3zcFc4DiNuT+kxPwFHAxqsM2JG1Jiw4a/04ccgp9F
Rtm7eSOmcHLxD+CUzlNGYZuVqh85FeWTA58AUpY6eDLH5y8TCX8E/kxVh+Mdp9+P1jjo7eynV724
WUnoMwnjqg3K6uFygx//wv0iTlhM9Qe1WODZ66Y7iI5CiqmzN9FudagVLAhgW2EwljhiiqOiI2R+
zIxYH08P3rqF4aeAGERG9TLOgUFVno1ZoUnrcsFbipExW7FUFgYgz9HzFlndISqDNlixfxhKI27B
0iL+VFYrhsfP4iCfv592zM1yYnVGGNVHu9jIdLkm73R4OxXi+U2b+DknMWQU2iPqn7CItfMqLsib
7s1Jz7LYVphFfAPFTtVMWAHFFwOBfdhcBWaFMvjeCKe1DUNmpoIhMp6BCeYCNlOuquNxZnkJTcCq
B1Fk0Pn/UL8wcpLzF+WtLq/zlIMcnX013W0RyVkZNNvF1hVVOf99yIEpo80jz77ijgU3aSVOrdGn
9a/Cu1A+r13ow3CABpG5S15F+a5vOPoqXbpYNl0TtamtRsmiW7l22eb3j99fr825QScZOiWyEdjW
nxJ5vT+zlD9qFN+MHW+lVlAA6LIU24lex4okRkw7PDT47i1Jk1S3/4RaAYjWr37jpdt8It2QRL4O
0SNfLAsbjTtGS5m+wz4vgLU42eeHT61wEKrq0lvxrLTSCHVSIwknvdGnSwKkbzpUyZqUDE7TLRku
Ztxs91ut9GYIW6emgn4SDartefnT8bEr3LmkozeEGWXWZhqsykm059SJR5uTA2qrGBLhgeMUROJv
ad6J/ZURcH1jDBVxMK9LrIcYrowvxVkv4sBCQAV0GwgUS0+La1FsQBkQxtmP9g6/ihMWHLeNN7K0
LtJLq8bLEmyA2sUgi34SR/ZDjiHp2YSKb+ekjnTmw8SprmMKW1ltuF2lfgZXm+j6bTYQ+CHQ/Q/j
RokHYKtqSYm1k+zNKbtFo27lCXHE4dDpaFgY7JgrDmcbrvVyRzc8hdMAg/Dxv9YTEQ3lRZHhO5Jr
RrpqczNDdof/vXqr0jPBANEohl8ml4IdFFjMlgLXaL8XOsIUThd2JG+9XkdJfmIVNpdzb7hdHBXQ
WS88qpRi0sIaQiIYrebl+PvUM26wkAUmrf3HdOWPtzinJhxD5BLz0Wt+CxWjENx1b37x6+XRKmwz
+BRCgIaLGGLYuEixfyYnFuK55Hf6mWKRGMudtsInxV7a2ptRhxFcOcphp5Y1nsDPDrGxe12UYERe
1tv4sFjf0BkHyosWQAOXTwE3iEPtuUoqLcwvwCQcXUKR2SkHXV4/J06OBZgKofYD5hIRM+p8OdqY
F5v3ecNIE86XeupluF7EwKQf5nyB94nEV2zZqlxJ0xwkbyov9b1LN76h8qyxv3Rfyd6lklRZlqIp
mZHPHkXkb94j0zTwgCrbZ1azVmu79kHLuvbkxiE9LUU5GcFg3/RBX8DTcjCxQe4oMkBXV+ENGqQJ
K8Y8UvAH04d6AP9Ai+kTMAH+D3G2pRcjlAUhCaTsF+HGinU4Gd917QEeWwlW+8TIWagVaAcKj//k
fqFvzfELGLJGciCVGCqq8+etuso00uBcic96QyF1UO0mN/48COpWEIV0y5/w0P+mX/SY09BV7RaO
CV42q4FPTsURGU+uEXCEnLgY/cSgTBjgHsqIiNUFVAr7yfIblgMj1uuOkkvOfEka2sO9MAeFernO
PBg9U4tEF7II3LP/QpOU+tlASuaYHClExf4qfJuoSjBoPLsmDoFjWxN7Wt63EqLvGXAHVaeSxNlE
OfeKKJLThRThaRn3E8dDKMHYqug4YqkDzi24WeMVV9gXWB8jXtst9tsvICnjEtPfU3iCMTigoIn1
jjkIKjF1iU18qnFJ3Lue99EWlbr2FbKXgoAyqPQzxeUqX1YPDFw+VR0wFatsUUT62jbbzDOXPmEd
PwPdg/voenhUKtu1czjH0WvxOAQPygshrX4TnzntQfiL70Jb6fTduXR5v30oqEdBfseJqLf9iKcV
fHcTshhGhGlY7xq6BB4PZF2v5OpHd+kUx9Xt/tLy2PQGbpfXZtxN5E1l591MpWxJHhxjK/Y2aR/N
V4hW0WCvVxcg5QfREFQNB/zrHAx474zJm9Iw/p4i6vQ87xV5QKunA/jOcx+4VmgkPf4ESCnMCEFO
pYAIvL+eABUrTq/RFAEvvMEQ2/naM5tYk/AK62PgsgJTtA1exGvPUlYuObisyFeq9amiq7ZLyCc/
6iw5cyhCcqJfakXUdd1NLo/K3ij8QNG5Q7kn7u76F6daXaM6yFarFVRqaIZ7UzGXRqh8mg/LPtp8
oZRi1up5ZGDCqPFd7YWUvTm6v1RZ4al3EMhMxZowJ09ffTyQY+EvecrZjUX/3O1VXbY1OJChtbI2
o7w2WyF6VAcFBJq1CnYDhbkkxbZgMAMXnvF7kGySj9KVWIroHnyLK2b9e9RPxFW6Ta6BhmUCdirM
mTTf/OHxuAy7MF9B+fGYNXgfAivxdgKgpcsaEy2SuiZghj4xENnQ5M4K70rLmAmPIrezObyJcPW6
pRc7dUGAOeYhCdl3eYxHl1jBgD/idrzV9CD9I5Jogyygox3alPE/u3tJPwF/Y2hK1/IS0zClZxIj
zL/i7tS93xdJNzlZtIAiw7h1s9zO0jcDBRX5IV48mVhYjagfHtxakb/yLfH6O/w1FvuBDZhvq34H
5IAnlkC6BVf1pbUMaa47yhMgEJFEImNBIyhkBYZf3uKgyW9pKW89lz+IEoUbYnNbbLUf/2mbhoF4
HnE0LqE3GoK0bi4x6mVECz1BOru0JHaOBXjO8HdHvzv7wQFMNmgMhSa6jteKDA1+qbvaWjgSiAbm
xn49RZL08Nrp7+DQ+9lRsChg9TLGsEDnMfBnldbY7r54XB9GunjcEJysFv0dXnDuMxt8/6guEDT1
S8qWOT+MpDvbUjLxC+gTWRQffIaOd8vJrP7kSz4BWQgjQ7pT7UGC+YzCl6YSA73Vq0g4tGzsFSM1
g1PKHuUEgKn1x13o41mtTzmy472aNFYSgTXk8h5+zrMMeU8FsRfYByRvMIvJIkGkKpX/SWi77JS7
sa1kbjXwdm66zyI+ksQ+oqf3bhdnMZRdLp0oX7GMuymw6oqDDUeT14NFolcoOMPkbiS5vsPj71DR
hjEpiUZhB/BPEYDgOnHqkXmEQCKS8oDacCG9VG75ro22tUVfq6C90+sjgjtMoKWJHI3RprD/hPiJ
PlJaHPbg1n+F8vQ67aXJz8DiJojnR+22XoCFzGTAmQb9c9RIzKMpmc/hUVq6SXCYJ7uLf6k90UH+
DGYUDW49jr8XSkPpNbX2DDWRCMmgcMz7TJTESFr+qqS7reX77igstOzpB6WJmIKOi80ntqoy96VD
hFcgxaogyXzNjkR2m5CN7ZQOYHgLltwC+LeSc4QW3xik22hewRkWKmbnJKQg/H0bta9YsawyRoqQ
KcQdG9Lj/A1omCC0uGMch/Br8ZOY+B1fzLRdhovgoGcD535ZHA6em5268W/kW4AiNQRnwKGBFUAK
KlYurY+h+jGG0Z9+44AXgZfFpPtuQ/uwTRhwQtA75ybX4vdIrEQX5GOFp9AlqdHYfoe/iWXkXnlw
Lx6QyxSlY8ReX7/h+STy9xPK4e4Frc7cRwC/3hwYyMLwvOFeCLj8BpmLWS5AGVzDyRmEM/ME7s20
v2/fPBRnzfbukcjdZvm6A0Ry3fmbauZ5rkT4cOg/GUPOjNh26j/mKdwoD7MJw7yUriYvysb65SF+
fGRrkUsczWj7EjqZxFmKSF3PbnIHeVL9Ygm6UfegFqF2UltWt+JWMYz51iDG6hgdzmd5HpPU/DlK
nQfILBRk/iaD/1W4mPW5bt/dA+uQSHQRXCpwW7AomOUYcVfOwch23A5EvH/2vhYvZiCOA2LXTh/I
kqAqWfhe8aebbxtNviP3rNety5wR68dyGyK4YFLctcQzKJT0UYR9SuZoscLl+FYoCD/GqQd+BqbD
o8OKfrdpu2+YPIqSm72EGw8GXo2UqN7lDW/rkubKcEoO02umqdm1sq0W3rWU4WxgmTfQdvbtrTtC
3ZtCmn+U8w/EJeN4xOuxEUZC48IP3EaMtjrnACci/1+XtWQm0xf2EfmUccGutIpTZR1DANuMcLGm
XZeW6UK2nIp6VY2TxpsN0VSmVnkGJ/jLiHFc1DaslugJg5inVHtTejKn5WScvzZp+jkXvF/a/m2V
kemyVXri3a78CeECtmHlt8mpbEpQgB3vv9ZJAHochYMzx6dgwxQeyey1TRbrWsl8FZVli+POKUvk
aNqgB4VPU23JwiEJ0LTyvtB57T+e8i8o2yKbhDl/V6TKeAGUFLaArL1BKmxldUkiqfMF3PBw7SKQ
xiuNFF33oUL3XAOY2SUkzi1K1Qn85h3IWElSpIGebd9emLk1keeuKJ+t1IYba4atzw87H2LmBPHn
iYV/6JaMA5IYxaDtulmXunbGKbYUmOUYkoWm4bOVFe/QO8XIB64vjg05BwP3fAj8m6UP6TSLO/D0
gFpTPk14Xedus5HnmZ9oM4U+oCoaQoRbI31uFIDl8V44vGCOBTJm+zXJLSAt192dO1B36WsmK9Av
AcxGrw7ZnLz0jwJKMyW0UJW9jR1tDZhsauEH5oI93A2/4Z4yKNNKYxh1UHT8pNiI9Jt3YCXkt9RU
gOr1nBoktFYo/DccXvZ36x4oC5eUD3pp4dWVeen1EO3fn1aOdYpMNA5JdbJwHd77Tj+tFEqK1wkv
G3Z6Ff0BFq3CtGTdxyU10RxenI6HM/pDL0O6xaK38nniyIm5H8W9mE/H0WWKDvm3ffKLQQOdHdUx
T8lCdOoCg0YTswF+FZ+wlxbuTq9mtMHB/ZCCm5SklOoxoja1ZDFOn7CUrySS5FA+OnQAJSZPPv4m
eZR3XWwMbhR0pAHSq5wBxH2brVq7TN8Krsk5QTpGLzWD5dagBSfzalLglk2gMj64UCkroEtyCiF+
h4FLvzxMEFmewhPOY29usD2nWURwFKTIeHvIhPRXoirRDzbwmDNMnQcbus1mP1gTfZa0f7lAK1iE
L/GB6HYE4vJDCCQZg0evkDueOCqI3eO+HtaKK5gIURuwo57ooYCU0SMHsMPStthRBmf1VDEAB6I6
g1PizMisHIQTII2LeEQcnkOnfpbA7wkenugnIr0+fO00dvmWnDtanu0WnAia7xpcDwYIOiaxJFV+
4T9VS0JuXy2QUA5Gk4fMtY2Z2BWgsYUjS97X/GcrVgqzSRszjb/0ZTgc75t5FG9sBK9D+lvKbBYw
NMysW9ENDk6hpVY0Ux297hofsXoWBpOATE9HTJg8aVldWqjwL3Pd5dc0j67dqUil6WxAhIT9RTDp
OBDFNcG5VY/7lIOnrwx27kK+fK/2BPvGCsdrVJNKuqrsEoTTBDj8vqXei7kM6gPrFkoIPJpIjlls
YrU6dgdXyx3EO9chONTCUlCyfQWG3gYkfXRouA3jVFMXaLCULth32DX4zMJwXZWf3JrYTdATEzvW
OnbBZBooqXpr6IQKw5SWHiRFQ3EU+ICCUoup4+L230Kr4Ua4dpb3ZrA8AkH0h3GJgs+XpbJ9hjTh
D0jMcqaTwobQoDLjV1uNMGa4sFEOObAQ2gJrlXVyZpkykPkJ3vcA50Z3UJ0Ki/5lUZirFeMmSLZw
WRoeQ9Z3IrGsm958Pv0RNhN2TZd9SgzmYYh/a5mBtC8bHazNnf/PeLh+7u5tA80uGUyy9fPlSNnh
3j8Ah9rJHRIl3NvGpgeX8n1H3kf6lXupZATweiOrBuN1Y3D5di2XC7XA+UToSHxRIm8G3hZWgSWv
aWADutpILD9pC0bnXN3NbCdjSy+v1mTYTdzpkC2SvIwH/dyZl1O4pl6V2PzXNa9t2qj2vb4w6RQ/
P2JHfJgZJ3OuKZQVTEojG/JbGcivgyeP1GmCq2gtMipJl/G4uvAhgtVsgW8RCSQ8CQPpAOyxv5KA
HfTbzdcb3Nn1H3tulGhb72js8QC/nnIm7/g3pcLAXoEA3nBu7LbZYjC4v0KlJKoC7SXQO0Ol1m+8
0BKZnDoZeuFFBaFviTWFeySA7O8NWedTnJoEpY43ghhxSQSUEs6ryV+stY1k0yO9YxVQ1dWEMBts
lbX4Gj/kINL4GOhLFlsXWJetlsSSzBjysAYlXyJcdONVDMa5tQ1Ib6/GEVD3jt3auwxnDs4xaEjA
lpGAGwlNjsBxP6KNHYxQQfOt7xoPikSmCwyHgUo8lbu5EfSPxfYqG1GWiWFjHLCUUqW988fZNmaV
g+deJtBSZQXMUxqQDrjisqAs8NZAiRBp6ADb9m0Jkj3ope1wVGixGe3DLGmI2daCuXtQjOER+SUe
cDNjLoi0oZlTWnw01g5HATVSG59H5X+8nMKjnXbGenhs6pcj31y4SHm4G113atnZrxsI/z3k9Chi
SXOhpRd8FidhC6WpZDMisoExd8G9xBPOYAtoDunCXMrscmq6Eb+Ej3gvdAZaKEbmAECPGycTUmx3
AA+61j/T0MG8BuF3rLwekmJ8OXhIrDRNoI71A1ParpXm+qAxlv/Rxg+sv+/K08zYrvSQZzdPILJW
qdTEsZQ4QWlKiVYHZLp6UrYiPHhB8trvOmAu74V4GR/LH6Ow5Z0cq5950ojTdWop3/RSfMbg9Vg6
GOBdhM4fZb63dI4RR6nWyljHr+ISO7C9SBBwKFURQd1FEY9jRVs3Fyeco350qzb6svgJiqxwaJXl
mSvUhu2dnNA7SQjoYZG+dGu4Qd30tCJbhMez60acdysKyw+cfBNtoBrzNArV0jxkuDrZJpNGbDVX
/25L/2CXxTA0n/mv2iIWPjn0Vcx/fVfJmDBy57/pXGKWDWWgU4KZuy3g3pP53uoDF5dluGMbsesZ
uVb7Zht4k0G90UrwhS24+SEnJlMfifkXXoeIigdjvCTiQiJ1xSlYm6+MKzMPIBMrRsNWtDpTiNqB
J9U+OvtAedpxXt3ypjlgFXvT4h4shAzAtv9Z+tC60cQkL4aKD993nXjmCpByEAo6pQpAPbNBuRxO
bl694imUbBPouAeU+ALYEw0Z2Bt+EviJ7x6JjIBGvDh/lAAO6uTxip+SObDKFOFhME6jrdDGPIFy
zNAO61yg7T69ytqNjy9TwEOrisCN451aAUXIsdOnQSBzu/R1jsn1fxxqtCtVY3ltYQz/N3CmapEa
ncKNY4R4sd4gUq3vel66LMEUQ1m2z3T1bKcYvAncwhoOmVkWE2o+BlmjMluiRqxh4abYHITtprWG
U6GSde+OXBFj6ub1CQ8Ng2T5wSkIk6GeQrDP2wDSMHQjWvD3SR1jw8NaxKU99G8bJgdR9zd37OFC
Gc25AuCJIZckX/5qI3/QXZB8dxFAQXkFxaiCL2+gSyi73fYp73Q7o7b7r3jCJsTRdkzF3rqGVgkj
FXxcCkT0/npm1RQ7BdeWUHFcxMUGWVBfvQI7oyr2trGV16cHob7tadLhFgpWDOXT2C0nJQsC4AV8
drEfPxJRxSndD9VcP5szwHspet86Rf4EORI/V6cFNGmKq2jTug6NuP4DiTleA5pgjA1pHCXqOjep
M3+bbKYwrL/8NQRu5040MouGaOfHsl1K8ViyZbkR2oK1bcT7uo+7hb9nOEY+gnpPSfwjXJ6u2Kh5
u29eTFpkcPxmrIFz7S+0f73mooJXpi1gNVwKxG6L9WCJMUcLiVWhhD3SkjyQvPCRMW22Bl0WPQ9i
kN7d6axpWDKEtGhPghl7jE3JmbmIlckHq3WIPb8N+OI1rexlCNWxAQnrHcIQHwBWIDIJE5o57RLA
7hYmNCp6m75hIh3JMcxbAwrK7fOkNpp86+llvDs+t3L0OgVCcn/gfElxEHTSo+xLtT0w7u+VVdDi
v+V3q86AnZAu+E2jUtYPArefXzo8cK44EY9/A+ffeITs4PwP0Lc4lwtY/s92RUMb33S7WOx9LdYJ
F6GQF2X9TzqqnwGqUYQAWZ41xJWl6VLTx0fVLLUcPysVSFSSwHnq3FKd7JD7E7Z2jXLH0Emxjbzv
+xIUQX/xOvzJPJd5zf6T3V+qT78qccIAcaSHV2pXW9q7Xz53J8/iAlVZn4mdQStDhUdt3vK0SIW4
ZKrLbd3uOVbzPhtXuxAIiDk6PILG5jHHl8Dve+rpOSP9T4Ljsb5zr6WwwPtQLH5BlEihTvkv+bhd
NWEWnhsG3ENXWi5h7pLJE2hMeFORvktMGCKnKL/ZUa7o40sdO2EHxQvxrxrw+WToXJ20KHuq5sww
pQWsXF5JaG30vLKAZU5d60K+IK0tubiSxpxAw4D4ZiVRjnhHatxYB5+wU0F26RpYJLrpY4exQsi2
NlK6hNL/tOjxJdh5BvaRcXYG1Cji+D5D4A/2c5aAmxMUqvMSICmvNIxMczEXWdNEoZvwRSWfJCJ+
OulqJkNdjpton4OVIIgcVFUHccLK/rvLcHg7vdTqqdCczX9PM/WOhrLRhheTrNahu4fY1XPcVMqq
OCJXXDRcy5Srs6s2+rHyBi4nkzi7893Wxmj/9i6zQUoj1yXoHpys9ftmBxIXBbRoUra5bziwW4UL
Viz5mlVrA/Rdb8FIqxBNPSFkWsi94aLk3V05r5ZpCNw5VM3QqOcgWiZ1F222tkg8qGvbCK8neYpr
OUU5Z/KPtJVCAtbC+cW+8K0V/omY04yw5XzHQ2foPRs01K1YsB3trOKg0VgNMOqEkammNHuOsMnV
d1TN8M+eVUnIZYWpXwvDdkTZzXV6ZmFUEjavEIwOgulaaIveE57B6wNPc8xcRzvYMYkSpYWNpc2u
fs3ISKra5wzCe6s5pvU7sZZRgEMrTQW6vYmVz8pwy0k3EaBv1Ghp5ssJdpnZ0J4GDMOWr8o5uxM0
zdm9jvbfbErG98E4yiownHHFh1yU6Wd6Zic/zo+tjY4skvR47vMWGqkKPOx+B26wwp4RxQLOtU7T
FxfK14dcU/u5lGchKGUqMmWJzaDxTI7v2BOqyuKpb1UxwHFvUTZz3J7MpqSvguptLAna0OWSG8RQ
ygmOZy/MmXBl19TC6qldS4rxJKP/WqWfJh1guu/X9ZqNv4lJ35nZ/dsNMlgotRwfsDY3aVgnKlFb
njly0HjK0LqUVOmFTV2XTWNiuss761ih+69mIWdPxCytF+GMb23ERJY1+HGwxm6WBH7Ldhxp74Q1
nbmC9f/m+W+sLuoqqGkcBZILPNdHyCF5fK84LJtNZrDGCexqnS1sHJNEZ9HU+oE/dLV+5tJ7BYLI
og1ESt2iJG9fDzU6pXby2X0ObvlWTXD6zTVApu/SSmRwFP/xn/rkAyA62KVDx6YvPBZrrSSPsRta
DgOUbpiAoo55nZ5AxFMN96rlZYnCT4zyg0smnY/JsGfVKRnoSAsqMVVhLeKghCHexajlTq5vvnHP
bH6yNkj+kZlcWBXDmRtbgOXQkGXlal3WBXABlAQ5jFivUsdpkuoFfnAjG1r55NoGZx+2LelpXASL
UyW8e1yo1sy2kqTkIeTZ3IKvZTOzqDdIzQ/jsJ0lpyHhhWmiY+DqNHc8/delsuw+nfmn2FHrRwi0
3RetlZR2fwfcGSyr3BxgDNYvrSD7K1JaS7WZ0z9ony1GLk4eGLUXf/wlCKxjwzwKlq8L+LEkvIOW
VZRsGbi/foFR1Qswc83IM7x0iWmEhmzASR+eWBvMoNsXedtNpg5A8EsEdeJUmEigndNCBBwkVf54
NxI5RdA674OQ2794h5ry0I/jQnHUITsM8/fJMJT5ewFzm9/FHy3s17A3I/0QmQm+8Lab/bUOMr9o
3RcXjb+5tWnTscAbfa9eBMzSLVz4yJ4cQE0rUe8Nle+4LaXfSVFUVzSE3LKVs6wA/Utbpfmx3ZHg
J1vnnorvc47YGdwpzuFX1IEn5phsFKTRONQp9142MKFR81x46Wq8g2ndl4kZsIiSv8sj7rPmf9vw
SsKTxOjGYdjfGVkVnANLHFjsEWNitdTlxaA90rlRyV6qzfs8c+Xm8xoQnmGJpm86QzhDDxDvlpVi
z0BcMFMDzPepWI2oFgDIJfNW8pPclTUCHhtbyS9xjCTnNMftFPcl0Ryk5Fw2kyHvR+F0BmZuyh9X
MNrx9Sy5wcdlwgZB2VXr0FsY18Ri3UV3IdAyK2q5dOSSDcazhuLz/bAEtJUp4e4bxf3Cs0LlHpoD
iht6isuYW/FoqAueonJD/C1HmHakXWsG6pn9YpoInLZnN4s24xHRkKbV9dJxJHrZitaOQdY168IZ
mDog1vaUfVFNXw310Z1rkl7P+U2Ku/kwgo3wEpAf+1QLbPOYU19tt2/7JaJDUZBdiEpi2IIb0Vo5
Lf+f+L27eww84f8hitnA2VpdtrP68fytzmAwq25nI3O36F/ojpy8vRpnkeAoKXA3oGVACVDwzSB7
PyeQwmmzCQLixmAUkqwJecS5D+iuGnEMvu8HfrSHntowhkM22Wdnjbki1eFpZ2VACPelsBDLCDsJ
X5f/MLKdXEzmlCWbtX4EGHLLvG9fC1lZZw4n+2WX5wweqRjzjz3XACjRKNhn6iTE6mZSbfJ+HQaL
nXGRTWTIryUhimB517P2p9zU1k9B6dUqQMSa80kZF+M7cqAf6DhI049TcgFsSsNSvlvBkR8LjvQU
5Gwlovc6dS1wqIAsMTxchpvxLzCQdJ12g+t4l2beyUFlF7FLdBND5n5j575kh+3sG/5P3jqDkNed
Fc2GS+z6J72e/CO6X8CaHlGOjh4It7kvASmvV13vX/C2kfpVATYMz1+DWEb+0K7PLcPR7GkWjudP
tNskhoF+tzZmzyMze8uIrJvSIiDHrTNVnuCe19hFc6szo19vNgeXYTtYF4CHquF8Cme1g2xPRGht
jrBGLJtdugTt7HXd5wBkTBjxsDAwJSApZdTEUUDzfFeGbH7TZvMqr9aJ6qz/BVwI8l42Gac2gq7P
0DT8xMZSP2dy4RIx0lbUH5J5aKIj+0MNlKsWlawbilPtUaNJE/pOEcUMW3pzpnMpY9qISVjKUFUd
tn+rL98W4ziBMrgXsu4w/QtivTKMNihJhvqDP5Pjoq3ZORjziQkUQZoscakdHlGAGBsM1snpJxbm
rQ2YcU1C5fGPYTZLBLfnmDnY2qJM5MyvYB2Njaw3EVothadFdxZrb7xq5xtt2L4o7hjPGf+WOm6O
BXx8oS4fPoKm4/sVYmMQn+Jwv1IHA0LC1O8mURTRGriA4SNpjJDsyATjPxOBMPBglZ5qVZN6P0hW
kwewIRCpSQSIR/iDUgdzBsG6ipoxn+QYp9jsHuuCwKewp+AgFxXRfeaOG4iFsab4vp7SPeFq5hkF
3zNHRAjzueAP826lIjya8yWs9lnFufU5F/TkFgefU91w43YW7kg5kasx68R+KWN9ugxLFeC9cRQP
VtQzRbPPHqTbGwOv2xv0Gz+qE9q7jFTqbL1r1TG3iHebM7XCUph/Pdi5Npw133fqUcEO6SnAQ3Hm
wSQw3DvK6ZuPcwiD0kAT2EJbDUdthQdIlkYeP9W/8eOzOR12H78LZe28u57sDRscrzjLxI7MiYx7
zDGVU20JIuunN6UHar4Iu83retjYnBKI1xz9LfWSxNztWjfZLX64HE/C+iw4oXd5zVCtqjqkBL+C
84PTi4z9/r8ge4MTsvfEEWMXYGQqHL+VLfIfP2onV4Ths7S3fEiGNlUaiFhWvX0T5fWVenQzTyS2
NeoqvkrED9ZA9BmFB4C5HkQH/aOjGJbAnya1liOJRIW1tN8Vj8zbTe6+KQpFyOPAP9EiRnxcM3jK
H/gnIY+D3SeSfLd96kIEtRckrUV5bvX78m1vy5dMekcmbAUMcwr5MIyEnHGhxA6wMtMKBsfzehpC
Ctv16kd7hFUo0Xw3awj9/vqjqRUrFBy0kyQE0Uc8l/fLpYln6RpZzq3F3KVT4dgcGITUbC/BRluD
xTsVNnXw/sx33KDy/LPzwkc2bNf28sRHqoWzqhXv2wYts4uycFt1B2ejOxjYbEUmPCjjKOLzMivx
3idWGrwEVtk94EXm92Ki3m2oyVZj6+tbgBauB5a9M7XlaRjC6FwnnUHG9AYpW1gEUULJ2Z6wkaGO
aB1XB3B+EK/7MIFfVx6fWKSNjHrsJjbNJCkAnBAcfk6D//MQX1jYyZNy6GjkhlT1A6gOBqRe4W5D
FNKcne7ElhpvZj4ihikd2Itb/m2kc+KvG28BNtq5VTRxGNgzqmlQqKRbakySWF+PaGb7+WQvLfs5
06/M4S2OxGpvxeBmWZMLhxTlgrL4K0GlgtaIoe6HXK0sfhgkanDhbm0yIqD8qh4L8lmw4ltH5mBw
9PAsnZ4YJUqi0TnhIT5q+aJfNFxhB5wmKjbJW4ZjuFMia9Ohayo7Lglz/x6/9l/+jxZdG53xCj/P
f+G4w9zyI6d0v9tGU2kHSggoMHsyvKZQG1NeD8zgKWnBvY09ZxCGimtgRGVIiG7ijhX90L9tvSHw
1qBi4hPJBc+v8GFMJUYhgg+ewKyVJzDT9btXcd90BS1qCT7/FleIdhTjv0ZOMFSCbJWdc1q7qZzz
CNe35bueY+GLhJkw6Y5QfYfJjrkf6wTv4a6x+kvNNUnSB6pFtuOB210Iyd28K4dQA7CLTvlabSdJ
lb9p41rz+Q5fBQ48dSiy/TQu5O7JD8rxBMmu2ccw2ajZF+eZKBsIZCRdV3MesgHLB0NgrnN2Jt2I
Y6SMtNnoUP7g0nPzIVD5CcBQL8ADnEDU1Q2AsoOnrR1YhOMz9RDokp8kZ+pktksPaaSII4cG3Nm9
hwM8YpoIa9S/q0N+W+aejB/BhH0P7goIOTdxvZprNtm+iJdDY2Bmr/X5qdVSorIVhsb+1YpAgQEs
MoSTVjEkRbxURsvxKZul6dbMJV0DKrVdXATfV7b3VFKrROUlYTilBv83Hs9CQL74Rt+zCG8eaeTE
5OV/P46iZ3yUthLb9du0V3jMm17AgMEDUNFtoFJ1QOfamqYtbVCJ/0MI7TGIbp9gtRG9mGF9/mk7
PuVfLFKXCsFIYdTdmvOcP/G6yfK2sp9MPlgqSnz2NVOjlHIBR7hbyDNvah1LBYfCboHdwl5RIfdz
Rtr46fsCkFZO1BlSN71eWEZ3AG5Jmd+91ige6PvwhHrZmljeQC/mFMQHfebHFKYQLm8oZoMWCJEH
oxmSyC2XX+8mKrPuVzJrhKundvJKAxjUxo3FRET2smMghGAmJWY3Un05Kxl6UyNXwwUizbNSMIgm
buKvFIpuXRBQrc3TLqQ2Os1WSrkv39zWq5QSXWiscPukW0rwF8L9vMH9MmiKl1QkxJCxyPhpCRLB
Bu94E9OJAvGOzBoievK2lKGT9UJgo/sS6tmlNoIfaXzb4MqZA7y6Un8dh24rxfFz2ARFBNzzY+31
LKFcWo/hX14bXvxA8ZS5m1QTfKNqJkD+3q/Z/48aki67ZQGLeKFG6VCUeqV6EActaTI6uEKod/Tl
TmcJ9bMpDlXEBCbkoq77mkgQuyZx1qie6MA7uwybbos7vKW3h4PXPzSLFEaKHJDURstz0+BC3xX7
q0lOUiuedFngyV0Nlg5hnP8l6984iDV1k+8dPpcup+W9Sm/zVSPabqA/j4+3gclevsoNCX0MtHrR
EKxv27KvRgwXZmjeJO14pzI16xgR3o9r51fmoFjtWkA5IRwE5YwhXfCIdMIjVxCOqhaP6I1D5WPF
Z85dUeaqHaNP/nmNzD5ofY31T9BE7MTVZuNRzesjrzYAEGBwQ2JL9uHJaojiC2ReFFNs+DhG4Lss
JZiskk1DuXhNcqdrSiIm6gEXY9BgHs/nBSQiZDECJCppoeYX69qty7dVzO0DNBq2+to3SUtq6cYl
BbUG8bblnk4TtXDYXQT4YJpnuhzzhWtwnFUisq+Z2VPX66LfucsxGFVnbpA0kOeaShOBLZe9lrAr
Ylyoxt5OsqPP4UCmYVGSasBlU140vcrpRXpsz6BTZMfC3+mLS4RrguuMHhC1eO3jqK31TA2BjHR7
LeGdDYO2coUsjENGF08KOp1CGEtQcLqHpjzc+K/Rt6Y+5hQhLFPKzIwcwot7Jy6K4oc3UCRtO7Hq
tFN2wz42svmKeU3KanzzJNFAN4Rck7JLV/NlAqTjLOygvWjMwBwEEvNpD3yo3cvuYuKBFviUlitZ
wyY11VRz7yy6rIQ9estDftn3CeW+yqSmyau+5bfdUdJ5cXtDRNFFXpZ8rQTR/uP9+bFtq1EwcCS2
4nPK0Pynhp0nyF6CzNMe6eWZgq+3LWXw5qEZk5xrqE6zTmLjd+5+R7ksvqVPrkV2RBwfG+rh/Hsj
0MRbT7wxn+xfc2BafrOv7/FYdgHOaergmmOA2J+55ld7nvcSHxviY9cv04GMv2ikbJJfMAcZS51i
+m+CGXUdfc7tP88Kguj0yzwpRT+bgBGHmyIgM77KJnrc1TjJLMDEh0Qw2fl2wMQohzzvRDrqoLCY
qVbtP0k+oZdTWDm5l62jd7lbC/MK4nRuPUDEwExVfS2d2OY78otnlI429ONhpS52O28w1xv3SRZ4
H+4fn9HhB6C/ANoJBQwOiduS971NRn+ogaBs89k7n5FZlZch0fa1qcESrSMge/LImRVGlPJtoJjF
rTm433PtaVSht27dHIWyW+Wi41ZXLWPPH/yELRgbWabvbc0hNN67ikFdseQo4gALaYCOhkHPNiRE
ihQnEbzS92otpegriIoeJXvdJtROExkOnkzXNlr4PGcbpQMcZqBnNzgzVUCbTpt1Swm8zXRp5t+s
iQJ51k9UdHhwyiTTkQTXQiF94lEu8LRsNRYvQxE0DUIp23+TjMJ46Zp0K4jtQ7942KxFzhYEDncw
DAH4gRlEzaUH/8knbB/QB6W+HNZDz7VPQ4Gc2v0jqQi57wAsP6h49rA2t89gwdAyTTMDxaX0s0CH
d/FehDEjIzYtr2a08yjmTZuzVbGdZzFERCp2MSIHsoG39M06KYrXZetuCnEpEUWda5fd2Hr0j2iQ
wy5WMXbdCEGWB98Q+Qzl2Wx3HUGprhXDfZEZP1jqDU6+a1EyB3rY9PGDsgGVrf1/GMJFk64VEfy1
IQzmn+LQybmgQg/XXhJES/wP+fQfsvQDDqT8FkBcKUwIwhpMtozFgDE+xHV/22rkQIaKzuR6p1Fk
oZk8QHb82cdPT3ME50nI+TtARIjJ+whOdjv3H8yF42hUpwfOOJNt68dzlCjqIRb08gLtuTT7plcr
nLiq4V+qvlkCgy4Y8ZU3XNZ3/wHisMZoMs9yw8yVyRDn84jrPmrNa1Laa8eqtYFGVE76otzbgEJ5
Jh0ZR6NTzy1hpK+PpA4eTxS+G6fwMDqqpBDGDL+4fH0COx04xmc/OT5Ren99Y3txKtPqbPSd6zOX
aSMhJLsAqP2kYA4QvnK0R2k5/J14z1Hb6AWUX/1pxkoE0rFncm7M3wJFZuA1YwtawUmQv2iYaoPK
ezGVbDSToEjyFQZrfRGLDiRVM4Eyl081CNrq5mn2H9JvcOvFdODhxtpX/oIzQjXqxg/mCdteOaXl
TrYg5WC5x9wu3BjH+eytej31AjslSI/r4pqowotCiQcuhwmUkPgnp+mFPhMLGUIPrQhvzx3ZWoza
ZrUqlp+hCpbbRo7R7fx52Gyj94BMDn1NrbrXx69j5H46ld+r/dVHSOw6VPvc4mmOScB8l+wMwd/1
kW+ZMY3pG9DuImLaKCBtPVaBjTPWUnFn3cJVpxIqZbIia9eoEY3BtT62I9W5weFdQ+Q0o4C5aVmM
M4eQstsRquBhuTFhZw0oNPKJPPZJhD32y/VfyGfsMTmqk7PZhm+0xdx2b0ooClSafkonuTb5NCAD
mNd22AI9fGxNSdVtXJDFkqkbEw5seij3+depRNrxL73+TBdfkqGoUley80zSdqX7XTeulEsEquP1
lMW1ghsy5u0JA4GWK7h61ykLH0uxTrVCJcpzcLlcG3xSN5W7ItWeRgSlcF56TaKkuT2ILPBvyywm
nvvXzs5X748I0dTYMNj51LqEGbI/xaGdHAmE2eF3P3h3SgNjmRNgd+RGMV3Lv4gUWPPsdQ2WNpj6
mt/Zbno+7iTqUNp7bcbn1K1c78p4lj8Z3+Rpi2pfMsXAGDVMmDlYa+Vz6ZA/p7szexeFIXxkbF2Q
Xv9MdV+WTvlbxj5fQXrkol4Uqjeb/m+fsQYUB7232oly0atvjAuJzlwzVUWYvWVZLNOgAaBc/mDk
12Rn/UqFtV2I7Jhs5qc584OHu1tVH0/QYm6QPQ/qx/5P3Y0Ew9pmSMP4Xo2ilfsyYk2heBWhgtez
LhXs8xLAQZWOsbAGyAgzC9P1Yc+JUt0nPd4tMY8Gj6fUUugyLCNhP/w4o5QLYdnRhc4Jk1Bv7+24
qfyG6T2Snx1ZJ9D1wUh9R26zrEGBnHXnLYMahGIS67FJ1pDo9sNtLuh/WJ/IOM0qXorBMfALQ0qH
9aRL0Z61pYtL1LHKObtDUViKj6dTInu/8MxGyjN5W1C7+whB7sgdrPkCw0ZzJq2TcZdHwQ1VbSsx
V3796Nzk3MY2aQgVEreLGJkCpOOXQ242rus2Z16fbY15EJ/eccPx6DynzopYkCiqbFRVGQ28W8OU
gUZNPX6IHtY4N81fosXoGIlnvvXqT6bH6N9Hqt/v/JzyMQtANXL+BwtiKbgjE7WYTu01+oACRfnb
lZntCAy2TNsQuuepmzdcInADetf2KscKT2qJLW6qZSNvr/ogLpczJjvEDn9g16ciZTACLexuCUqB
dyq56n/cdden756o+OCL6CZSDOFI5E9L3O4j5KIHphsU5nRL/AsxCfXGRFL8B1BIGTqahAf96paO
mre57RRMdHsBVdW9axJF7mxIjgV71uAvYHdy8J8t1ZEbp0Ze5hMbEMwB8CpwnhV1y0MS5mjQPQvx
kwJU5I1j5pourn1FzY+L99N136Tx89d4ZLBjVXO38FcboYOr2bzL29a0K78tZ/Kh6c9s8UPQ5gWE
iOpWrr0OoT5NsVt5+cGbAj0r82GegO7nrQosjV9leR7+FLOl5/2vZmANaNN6cITQU4y5IrVoLRsf
9xQveJ/vuSfx3SluL+qbky8nOscVdIkdeV4mO1EWpLMoRA5LH4qaP/9u5o19X8inypknCSYHlLkD
Z2GmfiV3VhcS4SSoUU7rUGAxg0FtXuCxmc/l99RGXB5mRRrHd4kzoTSIPr0sECel7O4mLYiAbhbV
jU2jN14XfZweLMkX+jdRHpEGTLHCTVC20vk3kChk3vfcjkBk+CltLn81pNtBKjtAfdjIFqhNtKN2
f5u+jDOLu7ajEclgZWMFeE+R03yhmrphGYGVtjWHlTc7o1EYsbRTDAAzlwp0O9NB2/Tuo+qfNw6N
tKbzdn4mJA6ExoT7AfBMGjzMRy0dwyi1c+pYWuxAzJ6PgtmnAzBVRx0SimvhYglOC1YAEzu7hEJN
ZqkoP5iVkvuWLgxrrvPSCDEuVYS6+EL7QpYPP3xwPCD1cFUp+MoK/OvX120W9CA9hISuLsBjP1rs
5VTPuQQmswroDyl0Cv35aORDmFm4kpC5YOES7jA9eZUxDVtiV+jaQvlsIoU5uYdRRJf9wveIwQED
Qw42W3U+Woezym06o0CEluacYYG6XEMSQh35UxPe+kZ/Onk992uI2zad8WTaMyd68bNR8wKjQw+L
Z9E8OFNpTmabj5l+xrESMJS50GDaqex8Uh3ypE3JXcuQrM6JVnG4nxki7dEOHtj4nr+j8R1VAHpL
HCcZtNa3AA/+nZjhxWc78E6eckJpe9zYad54tFt3jKiATGwTNhmz6ytd2hOOzSgIpsTiCCxipOcs
KRkLPorKXjqcRKz07X+H/htN980fAQTwRiNnIxSP+OSvwrQSCx39A3vS05VLXnIra98mKp3ekUNt
7lH+c67CCUEmHmkUNPfzMjOy0DUNYBE+rEWmzCQQVrL0FwLxqQCHmfbK8YTdPwAC6GGnGqvV6N82
AlHfQMzeHoWSWAosEveZ3nepUFN1yuZq9IcS5yQjWSRD1+HX8Id2sM2bs5zZ9p/DWVc3bJPxCnDW
Tb6fqqY8lmvBL3wp60JkWPv5lWbz8Zw1iUs9f2ODbmMpAtpjrKZKdp3qI4bBZ0UFt84N1Oowx8j6
UozrnIF1CVkL0/acZOLpXwdJC2pL9oQ6REGkoRWYwzaY/Q+P0Go2ME6XJ6oJeO9K48b+XNO0L2CL
vmoCqVjFZKyU+/jYoAyY6EsS5PRXu2F9ddTtmPe4OKabhn/Y2Ccol77UXpMQ5f3cy3MUi2rRNEzq
DS0G16J57Wb1JbCKLXNV7IKO+s67bIK/p3+l3I/0JaRkmO0q7XA+LKfCX6KuiUacLOXrMBmkB4WX
F4ktY7l67RvB/BnOUqEB4OsQL2QWJLWziZE0MqUTl+GpkY8Xfu+dOz3orHT9/QU4bNdDLm0aLAba
GDKxPzTQT8HaYDSMDU808YV/kRfNJDyFF7jMaOZOIeh64iJdXUH0PHsAQgULoS68ymF76vRDN2CY
Tz90DoSzH2NXm5d0VeJ0ofKBY75EGi3KZ37jjEkZ+jW/froi0M4LEc/CjG2fpP1FvxEn/hi15PrD
i8yqiIgsE4zXcEmCW9+3ShuzF8KXl8zuAgzC7iHbmUihBdiYQmNFG3FkyQbhlg5o/cogGT2mevXG
kULjr+fI4J+sGRGNv42sYhvfgCSiSM2UVmg54mKZ56SWx2aYNSbsTUf0i780kiCF1azl28Tdtbem
/cyy+94vv2r+OvCAAQXIq6OxDNzRUUH7tRqkokbGMP+cp6fVxoQLV19tXUQ5XiX8G7ujeVw464Aq
cpuazVyVx24DqbsVn6l7P+U2OjUrVCqLwVEjXN+ILFHFmBCotZ37o7Jyg8d9c1/fjdSHF6tsEF/k
qlpbwKmOiEUYLoCbRFvuus+H5jDuAd5PiwByLrGYslqFBQ8c2HD1UtbHbun+r+D9TeCIzyFKsMHs
NmJLcsX/y6RaSjmHkLVz8BId97Fqk0ipht0sjgI9cF0SuMdFts/WSB4oUJcidOqEfM5z42wptGDk
1J0sPnkDajHDJ7R5euGS+pOiw+fVn5yvuEjQoAY0ubn2cj3aeaRVsfgxOCWUs6fp+PBg8iUKRdFu
+YxyDOXG4MwRlDJBB+OnVt/IkIQN0t6bQD/ykREP2apY/nEn05oIMFUbZj627kvLoU5cbsBGBdcq
KDHbuvVvXnU2NhFBNWAFPmEl2jqbh3gqSzAAdyFN7+y3Li0yrbAp5ynkE/4iOYbRrbpyLeY4/gGh
I0Ts2SUt3QoO6a9EBcjnlDRbhezBxLWDp7l40EbTtceYUgmkxLF2DgNfERdYvReZCRwUuIR4rPIl
iJlKwsywKykeq+LWKf87zShp0K/fKP6fEuZxZDp+YIdFfTCt3AZG5gTsrWXQkvHm/25F710ADCod
gl6IoMtMvfBKuNx0b03vxbQtYURY7A3y9ojeS1LyOIPrGBcby5fly3pdRi0iBas9uIZNI0sjpMTZ
tasD0nMwZTmYiPqbXpSBnPBJOc3JmODuuczWEPjcYhz/982aGLjvIWMAA585S44RBi3OPM31Z4lB
g8RAHQbH83kywwZJMqgjGKXR549C2bpJenlEyJY8ei+n3YjnQ0Xi4x9V6ajNnDZ/lTdhhf8G/AON
aP2hJR+3zB40HCyFmrWNwMMBOI9YjeiL0TcWqk896P8xQvwQ3lrxpajS/bG31JahvW+tdvtJW5m/
OuAr9bG3TEb5FOKBtzDRwZcwf4oopGViHYosIuUUxOJXSP8Xi2yfmaO4CTq1BYxCr+yvzK5UEThe
xFTh2S2ABHw56/PcjC7yqTNfZcTnvWOgzuacajpH0hv4kOo+4PvqiO0TpMlAZbD28akFW0zy9C9N
rtLnPCOzmmgXZac2ze2994wq/I0mmE5jVI0AWoSAiZL79FLIHgJlWBgC4Ky5AepXpEAI0tFnP855
TLSZ+RV9RnUWbenWJeVOmYdNq5OUR9a3MZT0/bUjBEZtnbHkD0mOR1F46ke65UDvZo5LH2uOEoqf
s1ewcaEah3BDnE3VMZhDDiEkmV6qfnKlZBzaJMmad6E7X86EuzJdrt2cmtFjjhrfxRtPOY419aCO
CGFCXOmjA1rHnOnvgynshrU1blLBLZz32Ht/j2gXplwTfyHTA84fgmng8qW90+DAyaXTIvwTVFs1
/eumriUkQLqCurYMhFph01L1p4eXjaV/yQIF+OoUbGgD0xkmHXtP3FgyDXmmUeJdmCggHF0e2Xxk
i0azRyv5InGHSmy5hOZ+R8GaM4SCsSYdffVqJpaoTmDIybHM+TcRL86PXovELvnq7B8PmkZhF330
MesgdlrYrlnwIC1tFRG3ND562qgkd9kwb029ezpsMxCulzrGWUjKSJJ19ilD/5VrgmlcCDMCrE3n
o4Lo90pJZnEqvg+FiNBgZZEJOF5oh80pdne3iW3ZZphUspw7ph34iDlEJN4vodsNqsdgY0G/hBe6
ZJ/cfQvulbIuQhSpnwlKIilpqZE4H8MV56K9B2WvEqkfajRTgtoFBeeaQoLXRgw5RCXBEvpPTlrL
rpe2OAhJiWVfssgMXD6ejue6Br1vXfpNGhn8QOv8FdSwWAHkIGhr9QUeR9rWg9+Y2aTYGwhZ8sXO
uoWCLyFkTB6UoBhJYLRlltoJot4p8YHdVpaPG9jDEccW8bnfJ1LMWHQ7moObGcrxaziX5oZc6+DT
5dYUtjIbc4B3TBuKCgxGfPWTsZ/8dIOC+kqbezs42/QAhxrRYdevD5gos+2wtkWiWxcs84UxdH6y
hmzLpgC1/5MrO5c1TBORnMrrefu60/CK9+Aa1FVN7hlh4uUwDlw7/iBvWO9OEt7azKL7D+a5i/8k
LE6meYe4T0EF0jast33UQv1PStgWTaHnUNrmRM8NpSu1cXU7dkCW3i7HQswfm7gRl2HQHG1fE0MP
1mNZO2JjVMFKV8leloXQ8BgQZelNElF3GrEDEeA5BEkQUqSbYx89L3uxZNoCUos7oZSLG2uvWj59
IjL9i69nGlY9rW1pam5583mXE1ElKYQr4azibE3DzKDMXvZPxQGRmOpNyvnHau/WgnYRmi7XEaoS
MlQpsENDZAJbIAy4ndp/koc6dkvAy5PQfdcXBCdGNCMRdgGfze1C5CU/cNQHtEssdmbPc7uQjAbI
t040Ph+ZejPl++4/QZX2qy29Gf51+PwE2RK5+2znBserlhYzgwtjsg3Opvw9G1emqicUrrFurXBv
fwrLhNl3w0ilwzYjcM47rMurvLhxu+RWtAFqOd8OBmH9zWG88UEEz/T9e53olLyaWhIajHdmYZQJ
PxXkV0i1y1nmD8/PfmA/mkLPNwBExQNyUrPMMXx12TBDGlxHsLI/U5eQfFYozZOHWxyKyAAuDReT
7T82xn7yJHJeD1vXTiws/iJC05e55n2EFFmaccUIGB8oMlgZ6xXdoABHHd45uuQi+qz8KZgBDZI1
HhyNm25bxE6SY/evKdh8faekoslYJKJ/jrNN7LNWMoAybAyVaiuDdCTkCEJPHWQ3Ug/UKMC0Z/zr
G7zuM/mS6JUNONI2XNkv2DQ+3uC3ILU2T+iUVjIlv54kS2MIZEWd+2PZguRkSRQHBKloMNVjrQQD
XDfsVDNz1uc5SLoazn4Fn+2hZ1/t2JCKOHWYKuudg97ioBBvKPgKEWkAPnsooI10yhxye8xQgff6
HTTtGkQA0tuoIG8MCkf8QTmcZvrKYrVo28P6oZt6uyGYRgIq8lh7BiYq/ZBqQygrOwYRqLolZYSz
Bm2MbRGJLTOju5/5ZmDbM0EQckor41moLVrMXKpOZJfoPHw/5jy1ppUD8B+pwY7fturGV+Rv/kBC
yionCTp7NJIFXFdr35RxXf1ZsRATHD/SbHniFupsl04yHs75y1DQlEDA+4LMpENlV51ERorvmCuV
CdoJ/BMF7nifiyuh4tLvNG/tcieLCzo/opNv5rM/xcJxyfDcZu/JH9v4JhViLaDMETYmOJgwjCwL
KGVlidCVWFLOl/K9o9LLBf3P/v35MYf9lXL2xyQ0kSiS4RYV+8cu9TofytkhdUQ3PN02MXZm1rPw
+orwCUYOteD+UjvRgfpTz1IW5nZ7O2rJoRMk4BVy9yCkKM9rNgPwsTqqb1PYb2gbBR8RjV+jLXUP
tzUTztpQfbvuxcYhxDTiDVKAHIw1VdcQ2M3m4wbceBASAn1R87pf1bple5Jx9fpa4BmWt7XUahgr
84BJIGw7XyjrFPf2JRJAkGh40lMk5eam9LSo5jUS4sbbSo8GC6plchiyjKcQCPOX2I4eYD8k+bM5
ALwD99itsvkMacipD9SZJti5BABG8Bbm+uePCOn30Nkz3dU/IZM/mFHUdz5GXXalhZsnF/M4ZpBo
p8mhhU9RHYhIjIfKhpIHOyvZxoY8RGTDvvWfgsPV1ikgB8zABLYk+jKwEjfWufsLVN2s7XG2zCfO
GUsYCXOYAUMp1dD5LP/YLKikPgsl6hnI9Q5hTw+BuzwvNh7ztFPHOkuoksFvKHo15lxCbtLN5011
YgPF83FDcIEQWPnNNMeiOj1HYrgQr+csQd9b+YVuUPtp5tJfO8boMaCp9O+3tRQ6/pOxXakEGONT
HazKZrAIDmAl+OZwlww2kRLuWMBRfYtf0jwzd35T4Hn1GR+koMRg2QECizj8MXJxAa2m6fz8AbdN
SxIS/fDfPVlg4OY8GopnJfztag46stZjladJMGOiNvQhpS4CEeaKUfiEUYOEBGBchRPBiVKo8uXW
v/0dO7hvaYLPvqjEM0KBzsE7MSBc9vvJxC1Ga3/Ow8uzj3Mw+wM91pfMpRNnyIbJlI8cMTAO965s
fEltH527/H6kXzHwklyVgQe8ZvPUnpJcNy1NeZj8f7QveIymeYEoNp8NOTQgWbkO7e8sd3m9E2DJ
klp+XhiXbpL+E2MLYOw3duqiF9vspsY4i7BjuG41q+MWF6z4YwT4OUkrAW/528hm0bBPpanFF1M8
BwP6zGY/0n2at4jdPOxjcMQGSIEGBjs8tnVMfDkGnuoqYcTg8QCe6R/J7u6OYTyMf4r9yhIJS5Vq
eTYxiiiExYh2Sv9j+6Pk/WJ+ARyBpk/yFGCthWKs4dGWWOvwLb9ElVjaVDTfFKy8YDvGsff3WicN
A6Z5rsGUUGA77v54+HSBcFfLnnRmioTyVCRA2nm8bda0kDLEcmxNZxk2g6hxw1jz9vRp6Xy3/eTb
Ioztajm8xVNkyHwNKrDGO+H7xvfpPsbBgObIgqj5hbXqnFtXuTKsYEpQFQb2RjLsC5dSlTWdWdwK
TsdsntG7oh8XPHXG5wvi2iaUCAf5E5f83n7DTnIfICzy4sY2o+QvSTqf8axbzOcS/BmnCNh4a9E7
aJrIv2df+GgOijY2LLe8pQGs94vAAyTrCwTqMm0gWEE2boTB+BVSwtrCpYUT3QRTZb1hNTmF77i6
2stAzYke6nIqMC9lbMkxTh9LKaZO5hXOSfUgVZXqIyHFs7bxdw92QU31slWyzFdM55RcnlCBw4XV
60E4K+eIvFQiDz1JuYfykvWuMnIHs8ohqDyf4GnRkTihShoWC+yyHRjGt/10B9DrpMSVTkhFNoGu
0vbijERmyhnvjl0AFFM7Qr2lxR5d7n8cqHuP8kH1YcOOd0iOw68DlWSxUaveXw0JVLPyVH/ds0+C
VbuY48bUEqP0kIvCCv4GMzFQMsbN8cqLkjmHVfu3m9+N2e2lPglu1hiB0MfXgEOVfaDgQAlMrwvR
yKDEaPaEreo16Ixy2NVR21NAzXnqFAwaq+DJDOtM0/ndFOd98IVTp4njty3zDnDcS5qL5gdOue8K
hrpJeWkljxNrkeCAK3nlXysim7x9wmCVNWixANZajepTNXP+8LrE1AbJdvPJ/VElE/Qa/t/gbCa3
OZwX4hm3QYP37r9fFUrHHC6cNjbMXGk6gmu6Xrv8HYWtpxykHeo2yYVrrYh5dlKzQj0YwPXFGxOz
OVrvirkEdvcfmui+3ScrZb57w3pXGFyCFmpI3P1yCb6GEaOTU3X7BGjIsrDKSCEAHlaUjJCmUtvt
ccm/2fiQevZ3wkmZW0eF93A4AuTyJPh3gwO/4U0oed1XFYwWBlegSGqHwIiTJ3Q2I7YuxoPqovSv
jCBGcey6rmCLbrAGQGBjt+bmjEsou03cnElLrvi6cwI0QzHFOqWiRI0lsOpUXHDE3EoQK747toY4
I3roL0c7/ryuAnfRYCGf5+CONF5qjHQulO/n2teAJ9eN7MFmtsLgjI0wUM0CAAkLN4zHK/HQhs64
i/KslB+CnfJ4HRm9SoFFLQjvMywiPUHrp2ZRKM3K1pX58hXGqZT3akjuthvpOtPnmr++c7t7JGCt
k/QUX+vfilM/1c8ssHnVBFG755Yw748NMbeN17kTpkEy+H/z506a8NyHbntPq4VFLbOubVMwhCXY
6xFhop3cx82tg30TxCsCOS/t+1VHZb6BpD7Cq3Sa0kHauhNJ7z7EtvSK/R8oDWevJqxJk1v5jAG6
IByRenPduTHRCx8NJ6ZSgan4KKZ8pCCjul6SF3OgJNj2uqZCPeMsnJgBvs/OyEQCTspZiiMwjiVK
itvCoZ4Ag7oateo0lLlDoJn5y7uQkdSupg8vmJEfb1T5ZwWH10H6Ps4pGmJGvY4I80FImo8eHh2v
yy/9gkXIV7nMsFMDjvbunRuqEF6PfkdT/p90D23+HPmyNJA2iyDhARQL4Gmn0V/h9c1as9DYdRO8
SKFuksaIU3rXkDE0OQvzobVKYNokLgQv+e+yXG7q7SgrvL5JeCJuQjncf/oAQLysoNDzRF3Ju5kJ
cSQwhmpzlKvaDmEBR2T8H4LfOtbUqIw4ACSUesHBtEsCANlk7QD//3ojsW6VUyLsQW8payzD5jqR
3ocqeXP+EIijlHPHhsQZrEXtWrv07OykVf8KadIWOTt8J83Pft8v+qhLhOFaAICQ6REmcn98erv8
ONgOsu1ChiozkZa/vwl8ey0aY6SSjwriOM/p7QLP3BomRLdCxiSraPS8qBGMLxANSJL5mm+bUIaj
6LVphVM7p2iUSt4PTpQDTEF4rpRJxRhuiYcksuWmXt1yhWkIvwneviptXItvsj4Q71gYvleGliCz
FluDn0lXxUvW4sH8ef2bxtv6ognE9tPIwNYbP9bbgC28OJDwObwU++MXVAo8+MYgnQ+g91YaaveM
4uldo1FVHhqDZ3t01AhFdSMmRJ49JdzZ1UaAH+XBk8EQP0r9vLmZkqKuu8N3XgwEBp/lsdDfAwp3
ROCyYfgNA4msrNpF4JQEpoPE5XjZPy9LJZtGo3C6gljycpxNkwHiAJcfY/Zqjt94bohuT03kcChl
Bf0d25gx1ndR+XU3U/lDHT7ZV9QuNrHjGbHBhsQb0r0V2fpIBCPN9WOfCTBTagJeVJOnWoj+N9Bx
GYavchdpVwbPcOL/6noG/xDobdZaXHfIvmNy6G7xBTilmQZ8ozPjtdad63xYgFt7kyJxd3j6aGeM
bSvpoimeR7hQD54gnqvMX6UXJb6aLdHdNNHfKgS6GPfg/+rqHjE30wm3MLTeJikcaJYOnl0YaqLe
MWOwRohy+3gZZ8/sWHm+TqRP6N7Y/Tc/XLXkoysqWqICanWSKHdKA/7rv5dc4aSPlimp2J0IxGVB
pgM8lluBLgt9gqMqmdoTmjiLncHAkl1rnKJL40T2o5uSprnDnj+kZ5yPED9hnqW0WuJrzZpZl61L
AsZzgrdgT8U+Dvby2hNCV3IQYUjc6fV7S011KKlkFI+Z15K4GvdXvUCN7tGC++tNXTC2S1VlSPr6
irhykiYyFbjdWS1nW4FhEj2At9LvnH1Q4iPrOeAxbPtxWDHtwX6RVdjYaGd8qPhRgQYzoCP59mAU
h8if7N03AReBwwNteONdzglXKLS4uQUzjZr7wGmHM8r0jBBe+Q2EhkkHCVWEBJkdQueDE4tgACdD
eedUWtgspx2u4d0a368EneK/V+0yFoP9D5sD59ZAGYz3lBfjqgqz8kwzEVprY7sVE+8IDXwddAQr
8tOpDUomg6dbxFn/b2UfmUW1PkoLOZkvPLToJJMOGJS6CafLRn+Vzk3QzfPRaL90Uj7Sm3ShjvHe
Q08RSAmOz7vVGYIXYYdykdYPObONtU9rUjKfsJr7schMSq/n3DseygzwJC3Zy3NsCNIs0ea9y/M7
iPYZQnJmnv8KykLaWtDSOp1WswTvFoi1n/aYqQVmxd3goTp4rWM6mL2s5O6ZoFaZkStO2lYr6YZ2
VBywaoSCbPiyBxr+eCvzjKW6xHRt5PE4Wzh5YfCt2rOKtXsdzCSaRvTDiniC4+4phNNEoo/7o/rB
x+AT7TFCorN7lQyBfYDR8Pj/Usf9ytdySJ+HRbCouQmggakzsSfHT52QReh/wJk7/Bx6Pl2t604I
mFNMJ8q3U8ZS6fmm/0TEe0ovxiRQjMwojwFMnJxfFF5B9KdXF3rPVyMNc9R4Oh68IvIgscrBECg5
G1yJ10dXxzNRSg008mNmEmVMm3YobwDayS/xCdxrLTpVmxEfPcwsrF3gwSvmmFFqqahoF3sD2m0N
rOFPjHuXBQG7XtwE5wi1hV4xhyZT8Ii9pILqYQ7kKnEolMKm8WzZdvNi/E6Us2RIac+end1ukJhq
SzKsF0k6qnYS9EGseD1oMElGnGQKtb7e0dzsM8KZ+a++s2UrPZLXHlSKUtjwXdHsfouSitnfGmF0
z7k6dNmqOD/tJE09LOFsUyocRB550mBnBbsiFwImgR26YiqCW1Tttp1Rrt85sQeyehWb/0rrxvjb
36gjGz8ycVBpaSauOf2pIZD6fFtFBG+F+z5KtUraML+sHiioFQpM8uiKsbvECEXya7N3YHXkqhck
kHcX36/3pEbzqub5wf/AlcOWqWH2sHJ9fKy7HAKFCm6MCUsvp/OWTwsTttM2Gp1/iznhq51YAU9V
6eIBtebSZA7oYxXfO1RsT+8Ecn9P4aSn2puurg++3kG58ZLgQOWHQ4lrbdHMNZD6iHFp3bmyynRd
Cm06+N7YZN3dDZW52ZY+NGPpNZmMwnXk0rEIZrWieoLB39+o0M9jMAhOD/DUJY49lk4ddiuaVYcB
RILFAsUmSJ/U7Mk0AJ62Kqz1mtJBSd5nUTQBC4phmHgS9D/Al8gwXl8YjXDxKVVie/dOLOqamphe
A/y6YOrQ5XlSEp0ZfHCg+8uloMl3zIeyHpUZlbjYMmSCsiAKHysWtI1CHsONO5xCALHfV1pNc8KT
YIKCE7vryeb0NT86aYEVG9Ld91/OG4/VK7/JoyM/bYrG4m8h3M1H4SbkYWvdGNzL6RywcDdbmGRI
MTZIqE/p1NhFP6i5C+W9CJdrXMP6AdU0ITIDZnMlacSPqUT5XltmOCZG0rXbkhYbQ78FsoGQNA6p
KS/Ckvk/lMfzxrrt2DfYlWaJijKIWWdanBN6AQRflHqV+1VRg9EX9746Y/ocMotyUdb1FfU5drp/
5Yj723HSEXhBSxT/tGwdwvtommS4p8QyU1vKx4BWWmDF4beu/JClhfM5KTHUJjR7Vmmja0vglf0s
KtTaamdcEtOJG8ttQ0zxmEYCSjB6zt4zX9xbVcU/zKoWnhRjPyZCRpXwN0diF6A+YWcJR8DJSbeh
udr++fABeyMIZ++155SHZOiY/3mLGK4/LZCurd+n5I2TH5FczxvO10s8n6xkK9PEY6iE5eFc6GEy
AbOvvTsc3UxDziZkVCMtYTqE6ja/9dXchHdBESfanH0C7HjnGAceyKP33I8fuSabBbBJ2QMEECuF
/OHAQ4AqPsp/d6tDHU3VnNdTtlCQchSK2HA2RXFwFZImKlkKpPwA4dKjsYSm56JaQDWs7VNR3EyH
svQdFOBlCfu6mo0s4nwztoTngk/8A7s7yeFC06FLGrBEXMPaL4xnQeTZ8EG/zfUjXqGtG4r52ocj
QS/Cqdj9l4ZHuMopiQ6ylD88iNptq+LkcacW7vW+uryYPuSRD3c8UaQjrJeduQPJExSoodvRweTS
ifinwBVQs2bjnk5pztk1dtKCMzhlFIo5Fp2DNn0JPoTLWgB6yfnOjIcgzwwsPVCEa+cDKCIjjg24
DOfGQU1Pyd+WlrQhY9UnanARp7a5Cw6Kp6mQwA7IO202MKBnIQ+79uUk+DkkLjH1JYBF+RcrKcGf
GPnZAFa05T4cuYKuUyFATQrFfVAflAsBPW8a5m6a24ZpZqgntUgCCnwgRUryqEBXam6uRzK212af
K+OxoXXc9E0mu15rO2qn3B69oq7h6pq4sPkqH11EkPcyJ3Q6+TVd44nL70dbL7Cs7wf1SO2hzx3W
/IMBvpiZbaD3/x4Z7cX6z+J1ZvzgDfyB+SJhePN+HIsYj6r88i0QddnvtWR7B8SJ9HgBKmQR8p5M
/4IaJGfQB/nWrsQlgpw7442cNCn3nYuQzCHsjK5UBkyTrKLuF5Z2UsV6KwgnaBiZYmJierOwCp/Q
Ro1NXhOP4p7z6/HtxXLESdi4pKkOQZtCrhFCZvXtxTXbVJxgYz4l43MCkdcYdUMTVGXsp5uv6vr8
nfTAzuPJv53QNw86SSx6h6vW+sVjecEDBMHOIvzwzkRoD4pU9+Jd4w5PkuZHicujFI1KgKYQVBiI
zVKHL0AqlmOtPtDUiMtGhJqPMFNQniWBMNVe/7bBzaTD003Rmct9DTGcN65Fu+ri8x5WlruTsl7k
kOz6B/qPJAP6H0hFgWoVUKaXHZwutRt7WAsm8NMgH0JuKTsuRc0jXY9mkcNPMxCAFs6bXZiJlD2c
TONLS3iiap0AAD4i/KOtSBVPyYVjFn+lyVKThDP1Rj3mhI7HWkOKtltylYBo3CS1fCLR2r98p6a7
UB4QZjxSA6uIWlMLq2jnZbheEoOuPZa6cF0wiEub3R6kqzk6314Ql9H8ImpvCPCN41M4NgmBoWUy
3F+Qd/kmFNKfboE/qLxlKIuTQ44pqGOXJF5leYd9qi6XLTHZNEiddfzVVnGDl5pfRWvDExOWMLSm
oqEXdBbXPUquA9JMupuCe70OlLdLB7tiFv8+x6pwALw9i8kxAv19EHUCtbIvnKEusKlj6+xAblDd
l/3F+n2LFdeDbSZTniW2hNZhEq9oSLBbVkQDX5Nh0EJh6vbEt/SjERgqArIQAGVSOhkfWEwByWcm
Nz5PdwLTCPo2XFES+VSociIcWz/jkERTyGP0+m14yau4fVji9fZmSeDw+BXODorUjL5SluTkCv/t
KkUHu61zsN/oLBu1KEETvX7Lsp2HohRqtb4lAjg8hpv3SrItr8vybltCQpKV/JXkA5eRgCdsbZWb
wpMj3UwzDXFBx1B7gPEv9yxZb4E4I1DqTOr0AuqIXrC3eYoE+gUKbaCoZR/nCOZEvUNkCf/nSeBC
FB0wo984kQ3TNa9Jj1gbTbOw/8Q5ZkOoCx8ztrN6gora3euI7Viuoi77asEvSwNopXIuLcs8pG6X
7+KAfGadIwVyfOR8L5MIAdoU5XSpYIl5pBCrE2XSXVTlI3mStMolplnNRynTCepQk+Z0WdcFQQX0
HiS+YK8EsqKyYGfzhgNMGRTFdWd0hl9nP/sAzAF6Eqb4ls1ijs79s6H0gaSqveHXuq70I4WdESfo
zFqw0gPTheekbJlIVa7tjBrFzAE2H8MJsMEH8qU3mvVy/4OxYhGIyI6cO+A/nc+VdGTZDAu2RRs5
GfiB+VaRBWY9O2XKxIeaueDrFqqNdbjlOANHq3ohw4FjFpwJW14THeL0/EM6O+70tIBJHGMMYqao
aU250494jb7kDXbwyS19tCQizIw3YI080fnS4NvdOIUFgioz0IB7NW4SYSOXO7VXLgyx13LIFjpz
yYX55u/0HvmN3XDogrF6rqMGZBc74NPGHgoKiRlAiYhLDruZYITI6tcQSBByLtP4K7GZhLGi4vzg
2GCRXfObGrXDMvMuVjLEhxsBKgsenhyRPqY1xRJRibqtn++rcDxdqM/kfjtRdTUHtmMyqJKbw1cD
MMoAlh0OkJby3KdlmSVIX4MubA/+oQ4vhO4+fW/zGPqK2kahD6rq5nYqRBbJxqe4MWp4/Br6OJcu
PNfeGruofNMtuDrgrkU05lSQFCsInWOx7MqxvaeVF8cLcxjBAf2zXvS/KXDHOIqmfkat5uTfstfb
k4nxKxYpucDdWXFb49nln8uRWD9Y3ZdGiEJ5rmXQ41R53StiU46iFLpy/XDfxSGjMIooGJnBdL3Y
PqOBecoMkSBYHLb4MXxXyQu5NNp6/zD3X2BNKJWgaYMXIbo43cAQSnQHAbNad43kbbM4bCFylgw4
FxxH11Y6sBZQuGDcDEzxoSRMjeN0bF0jwZZo6HqSNEyPA2Cmg+Lh5RnAKQLUfvRV0lGiyNbZ6Qii
AXTjR7F+8mXZV/1vDGMmU3I4PSyRXYmVW50fym/zm+WnMu0JEB15FBT2k988AAlGGriUp6rRxY4N
YGrwoqfYS0/n714097utduEiRXCQ4mDV7qTOmVi/5gEd/ajM/6BmhOzuN+FSgSLGd7yAzCfrdyja
NAQIlVPPdugQVYLiubd5+9KljI8CCh8Iua76YAUzLU/4r2hQ2QWAuhtwRnjjGAQ3QDcL1wjP8XfU
KQUbhOqV9rByuQmDs+vtiozDYBb2yywu7Y+A/kX3Tnr5znZX2egPf2v1rhYOLzagahp8XAuU3Q/V
41fqOYNj4nCya+XMjY3/H/nd+cYg/oSF+Ldds1YOCkeoFhB/sTMmy/wC4y/TyF3iioD7DCEtu8iR
uzdAy0mhK8LOmhZ+f22J+WhUNx1b0XP/DTLcX3YmMl3vimCcaXVi2GrlA50iYL3L8fS0UskZE5Xu
7tuJu9AwITc1Jrp450Db4u7LnYKMqY1a04O/STBs/aMoWEXCx+MojBW3NyD24Kje0rZswE5SOEOn
ftl2Jz9W/WTZLBfvwrmJSDP5XA+QaxmmYq1fn9cRDKecwZqi/Tsf2TopczKenQNb6AIGY942M1dY
iAuMf1/kUxE3YbP9X++Rm36hbJtFrvwrL830BK0Guw4l84X/2wJ7A5Yf+hFEhegqRQGEw5G1B20L
R9+vcM2j1b4klif7S8+0yyV5EOZ+YSpYCVGCn4+LwmE/5CCZqhSmnCU/ReIJ8TJJ2A3aob2YNOBe
h+KdGsbzTdL0D1socEeOa4crP07rykq+4/Ss0yI5N0zP9qA+/VJ3SKSez33czTn7Zx/t9ryOTT2g
iQiQeyKnKS22+DtlqQNgoQDbfjAMzjA4Fili2OCYE3jq6l2lpKderClDPgXbT3hQYVe5w1N26mA6
15Xs9ZPwrQAPXSQ/T+U/PhB9QMptKFHl2E0tiYWQOBHyVj7jaG0mgpWULVPjwTVqwTA4oJF9pyM2
JdbJYYlfs/EY74eT5OQa3+rHFdSFRarx9hCbR2esDiYcMh47Mm7xYpeLADrqvS50l6WA1yRSwEZk
v21LSMPZqiOGUq8gT+THDEGUMWbggkk0Ffyli8tUOMqiHFCiDTbFyZbY4zDJSrkisNiO/DAhvN0B
wqVovfJhJtPU0QzgQ/I5FGg67MzBusLgXUlYT0kngpKdMCIQ9ER/kWeYWH1jgswpmMFS9HZx7ivL
IaP/zGXHON1k3qj7ukOyy/0WEWmwVdaROZAYhdu4rmW9UdMFozSQxc11yfprtFNU3cTqGfCARVas
Q9oVMBGA1Su/VCccWC0NUeuehhmuKzx4/P7m+g/MM8HUobGmmLcatxhNNQItNInFcEaFWeeRcho1
aWsiRRK0ncQzgZwB1yBehUhQh5LWbj4ubkX/es1ZRNtSG8y2MFrCH01nuP3BtPqqrzsQe2AqLCg4
2UePhOKUBipnuSPoBXrE2dsplW5Wm3b1IrLVR1ryVicSjBhxb7PIiiecU6Wzn1kWl0GpDzxsmEQJ
8Zbk8X/uEQOC1QUHAMVwvh7HvGggh3j92ffZ6aZ8Fgyae70E8EDpzsJP6n2UItKeglD5JIs/sG0v
S0LghEpSJ3vESiNb3J2DDRQbSEA1S5wvmcoo8AQhc6zmI5/D0X4S2uFnf7wJQYkE/o5nmPB9kgcs
+6ypWMrbiooyx00moCNqhOt6V11hBkC1eMD8YGQN7DjM+BAF3c1RzEjZvUfWaj2S3XCBJ19loRnH
z2pRh6iYy3S0NZNr2wx1fC2dm82gj9SPccdi/4LgnrSvT6FZvywowvNkJv89c+Hk2eX2Fpk7RF3e
UWUBPoW+emIE6+S3ulYJUrZKzJ9QWPQz/6RzpwfgCNja78pG4FNfW0YPlkfPeafvQPjXjnHW3BSM
g3Un+QC8SX4Gf1D40Y7sBJmlLxEDmPiRuKeL+QDZvBfrJK5AbztoNJ/h6xQc5OJygNrdEDf83MUZ
j7KcB8fSRhxJyynPHwEyQdm2O1ObN/0YVTsG7Z+YnSvmugLDKSYGok5QuMzlrnvot9TSmc+X0rOe
qcABFaJ43Hvl2M1jD+FpLKqjNz7vKhdaiuiRvSOjQm4ZWCCs6Rm4HIuTJ57x58LkplhVty2njT6o
02ACDsgbiq4Buto6D1frWt3Jhg2w2FFU03AyX+xKe4vBWwW76Ip+XqvVDP46+QWNDi820EMMWUQQ
f+fNfHR4mwzXWweKipWiRW+vWPg0RCNY69bnvSww7FagcLI2VrOn2OQSyRMsBQajKK0YlCrMWRQB
y/or7BIrZTPrVa8yN18vw+qFWtav8aGabdhZcXQVIHbzIUdJ6RPDvauRaxwanrX6zlMuUE4vPXsf
wfTJbLt7VQA+aw8BTrG052A9k7ZKDODCXICtLoQ558ZaVw/7ZB0g1Tjon2JmVKKG/Lty76+Pkc12
+7xxkzaxEfwbzOP0wpzMP0B3hxC+w/bJCEcQW9T3n3ecYpskTbialOAXWiqR1LAMTfLcL1JOr1eI
jd0IcPRph3CKNkGnS3OuzJgLD50l4y6CQeqOE58zy2QMt5GS+jzGfBFOjk0fuqFXRwoBflaF+v33
XeIBwFn0hRz+jyi96UAebupqiQbtn3Dl2FaxG50hyKPJ2pXgHbpSerq6KBvfwl1fThiGpvscCMnS
Fk8/TgkGa01TO65fzfPKZ+vFWPxJaA1DJZtw5u415/JWgcQ74elTqH+9cOuO6zeCjTAkV2aGw9My
n1I+EvAoLngwsA5fSrPTEOjuDv7/uDCRw7uh8st4j62Ib+Zfv6Y5d2SJ5P0cNFmEZmjY3a3/RMvW
3KYSr3+x4eqxgYrMh4IWB7GdrcF21whw8/slxXCyvKq/5cTumn+zlQPg5qdSlh3yvOwEt4Qf5N1h
5NDwHQNRIO5A7eM8MXuGGcO/74rRtzE35NzTW5Z5k7U7yHxxQ8x/OLYgot0k2k8SHDRzhuKLODdy
wr1hTRMrU5c/AMpcwh5sI4LASLWR/1Ul6VQQb4FJCd/ZpOzjforyVLtXiaD46ZdzJXTZ5kYtBJft
p/VR756b06IicB+plVMXCXlfwlLyk9IgqawNpUpK3mDtqs/jm6lZZP1Q+djDVvHzOt/UfmIwZuBG
Auvvs5YM5blCjkBsDNFX58I9iM8Bom4tV24kSD1nRfUuCuDsEkVIletOkaD8dMY3z5ldZESgv/2i
zRu5xWig+wVYK8yx2WOhGTqufP9ENBrxVp5WHidYHT/aP9HjDvJj0dytdJkcYXjIWjGfowsmawud
htXpeg0uEu/OkAQ4+NkC/N7bVbpAOflACx6RedbtLnBbkQ1QfvGlpl4aZ73bZNgQJ8AknwRwyt4L
T6Xp3/WH75hbHQ/xVAo7X8Z2ho5brJaqId2ncrMoR4Cm5O67yL9uYyy5uwzyDIFLZ4Qe9xEQ9o5i
ApOSoOdtJvBxHCABvX1XH2A4lzT9x8+koR56OC6YA0zywakS1jkp+IGQOpmN9Q6yAGltNlbwvw5j
5NdGSnjkg1wyND9VFuTFjhnROaF1jmIL2YMvfvGSJ4bvtVWIqIdEN449mw9wIzujTAjRlsdkMSbk
9937GW/l1Ndb1JA6hN071AaE3dV+mYPut8EDWjzWSMutomHzeXBVmmIpvmUPdVuc8U3JdQCe5qOB
+jmpnrtJ2gH2j/2ow6ENT3GRDjV0ufmxxCRFtg53GLXEiS4M/r6iWgoQaFINtycfwdBvlL+HPigB
6ghTpXtL4jPwPY+DwlVed4nbmeQi6uK96g+fpn+Waw2qjiTbWp9ZRqyI9wbPWLDZHI30Qc4zoQya
0F2gTsPRfatp8YwJU8fylwx5qlDL4FuaMgFBTjNiyrE8wy4EFubkGmPORc8ax7MgVtQ2wJhCE2Zi
oYyD5Z4NZY+8f9XabDcg8h3xTqjANMwSTFY5dFlj1PCzr5d+IbZTQPxqg1t4PSk47+qjWTGLqwp/
BhbScwy6DuOPevsgxWr0kDx0j9+4Ym/hBa0O8tLN3jvO8GoLLVoQnou1PkAmc67Pu0jshxCgKyIw
c4VZhhGzAMBmf39Huhb127usvJxX3JvuJfMLnsOtTRqM+YR2BtvBvwYuFTdUBmXR0t1rrH0lAaA2
frW9DcnlIc0//FgltnmhG0gnc9TH1hreBGRHm/vvr8cfRnOgg3EeBD15qEqkEgHPDMGVcJjoWR+U
5zVir8AZcrYpwB8GuaP4sxGSSFGwM+9nvlfG6LU+FNMdv4jASKUy8Ji0ttqIAk4tXK2myk0JfpUR
qcgz8xjXexQkiRMkmFwqmYlaNdCYmOP7ogNbpVJdw7SHxhwWsN5NDAwlX2baBb3cqSdUw0KzrTZD
QaZhhhd0s3MW8t78pV+Pqj9hqNchjPqG/uOxEDFGpKKsz+lqU+JoG3SsVEPrFGFjkAO73p65YBRr
S1MJ4G0A+m9jIXnX7U2zD9xjmJe0O1niAZGXFbG79HFQ2kXxUwptKN74m1NSqnDyvvKsYiwPc/cp
ZQlZfcJDbe1yRINzccam9pownvOfK3BRV2g7Vsyq1ZVn3vgZ6cT/YkYDTUcciIWmCyyKrDs9GtpN
wPH2fV8PCeVVCA8oRuBiMvjiIecLBbIjD3bQDPbKT/FM8Cr4jn8/N+ydRYWSPqtkbipMjX4DRtX1
FbYqn6xqyoz5TgxKfYgkb6REyzC1YfNyGQg40lE6yxPfX28B81GPMiTwPF3exJUHJgteeKkQd72F
CzwolLH2kRxCx6xUQ7jHDXxvRF3Su5p2ulWwyxPQvH4XqrLhGXwydqMkp8N8fsASGiQ/JN7P8Cw1
voMUSKLEBbo2Sxhu+s41QPJin3oq/JvCEXGeT0lV/8LIG7aUaGiyQFe5X6zcojNfmSfyKJYykHCb
1bM0QHK6SByh5tLKMpN+5ngIGm6TJursdxok7eAA/KkTQaBE/Sg9QvbRYvRa2PIQuj+gtiAojR1D
fVanPHt9MVEyBIV8dRFIUy28ghZc+lYnyXLv9/MwBEKAgJ1gl6GNMJJkYIPmS9ViIzvomF6mwlLk
WZZu+3AVbONk25kDPEtK40psAQ0UpfvSD6Tve3ANeBqNTSd8hbZk0mZ8flDNJK2TEDtTVpYaoMQ9
Cwnwwg1RYbdVc3HOlQxL9R3Md54UyNX/HkYtHS6/Dlu7AhzRrqucQau+CC/GSUkMXsHFU/irRN1m
e2bh97pRP+3yp4jlAZRADCGXzDAEaQo1qHWXp7sGqmItL8TbBU1We2skdFPP4HUxdK6BU+EC5nvC
wH4i/gfD0GmtRqHD6BbF/F7PkYNV3A/JdvQ/huHsSJfQaGq3ZwJvPOkm0jyzcfeu6ETrkiQUMQCd
LVyLesKOWcegCMzkwTLNYNfIgEpWljs3B7HQ8+bcYzQfp76TN25UyETb67q93U5kBmtaL8IiJRxY
RmUzvCfIGZh9uohEJIqkqUb+b3Wlg/eKdm5oAuCg+5+vHv2xZcl6FQL9wA4n31klOSFeR17/NHOA
LYVvW4oUIKWLxNGM8nJfOXQN454SOidjVgnvVMhUjJx5uoMn0modmd3yN6UQ1ivFG4aUw5Mgv9zI
necqUG3pqphYUbVX42tN6a8irv5gAyO8lsSwKKdpg/JgeT+XzHFJ6G8ui0yaPwoFrOm/Ea6kPeTC
sKEAQ8FJJk6bjRuy8/DYBepXsINHC0TZb1hIRgwOEKvxdLtGjT1bIKhAtta+hWhqMr/JKFLi9EAU
+OfkNebdUvGqhTwhaYZsD3jtTqxraJtE4oUMVI0GNALBuC/nAQl8KC8DbzBjjC784OTf2jZbj3YD
X5CoGrt88otoWDeIJZ7wfHfaHhzvCCNIXzZmHBImHbBwkANIM4vaFDsshze2WTUn/uCogkCkdK9h
l9VjrAMrynY4Lc40d835FcPrr8FZo9IsO83d6DaHvNroGaM1pqnP/+tDM3ZVfch0GNtWWOR7FRDg
kA82nYMshdSW+aQ98Tv/3oRCL8o1VAWz5O25ODA71Lq9v83JYkS5VeSNYN1SPCrSTyZgaatyj7m0
XNukj+l86psA6Qc52RdDiV4wiVf3k+rodvY3H6NfNTbKJyE/8Iasv/cbMsLZmsgX7brRrLv/+dBb
n6xYtzagk8TyuJKj/oh9NSTZMLrU/Ujvwj148BE6tm5VmoCtn8tiq6MifaVf8NOGfG1K2d2Youb1
tB+zvOrimDpN3RZJt4bvJTZaSTAZPjvP4eljPdoaeGOX97osm87SWcKn7NLKItI7bM9YXX2ikYWC
c8gpuGcU8so41vbHobNb33X6vCg5cMc/JznfJjzITHLyihoYyTEyPuPmgfiIhDmLEBkStgneyY2g
mgyHC4kfjYFilpoBKzFwMxHsXgAQJc3G4yB+tl+ILNYcUtt+ZsMwJwsA5tIo79C3TTHG18IOLA1B
G+37N0kMDuGo//K29GjhZRnUt5r9QXUIAwVpCZkj/G3iWs2P9mQByHW0X2pAlp3dXmtg35UQvtBB
PhP+pcfqQsdMX6sjcPCsZuZnLAcPaUFUm3YX/CqJJzb8nKgpLe85x8GmkifPHgpqHWm+F66H6Zct
dR942pVcPeXHX3a5qngxSWLWQ+O2l0x0IgcdaghmUlcIKHkccoEZYedKCZMyH52UBAnekTXFtYJJ
2Nuov4geaQEpgKb5gdAqwfOz/AXBw/AiB0YV3hlsL5kQkgt4VQbURvB2mXt/+KXbU2g5eJnjHq6D
DLVDut3cMLmqpueFL4gVNCgU855M3kPOCig7Q1i4C0DJ7N1v2eIyFA/B5QqUfub8loC2o/8g3O2R
+g6Hx/NEBVU4Lvw6IGUPt11bkcvkWFjyklQDcEaI08bkIHsXvn5BazL2sdud823E4UHWmhW/ER2H
pfy7H2fDBgNgWSqoWJFPxGKwwECM2TghYJLioSAfbH6pdatqyFcYakBGQ0+H0/12jWSfT99TUcEx
S6pPcN8+ayV3nTJcGEH2btMv9dAi3DeYbILokvXAeA/J+1r+RyWBVu7f5E11ERRV2rnDpzYBknfg
IZU0xDLWLMDCNUFLYBXTlJuCOABJl+HhDSlZ/bRYSN1pXeAnKZXEz9WkQ3Ai/wrMhap4EnbN3e4W
qjmji+DEpYqqyrxpra8xHzb2ocAldx3KiH4ovL14lIbSlg/F0lcVIHNyLfcAhu/eeOP5g0r/hPYs
VM8MiSQnk7tw8dZ8s5ufx42P/6+vm8UGXjFpfrCaSy0Cphv0CEpSfk3PXqZXdnEhC6RKTb04Ejb4
K5+31uqlXbFG52OiYMv+2dts9SG7FbjRAQDJv9+nuRi16UOLS6jvLPTE6nfhgQXsWrCZFnooPtHg
u9OpPzyt2ptZOcSqBj5b7FeIanoWziWfClClybZuyW4mzdqdPw0lh4QNaofxmosOHVhrN0Va4X/Z
okwVqrrhLbyFKlBNLArNVkH8ult8DrcGZVXKeSfUKPoD7WWjzh0Xzps1EdV51v0JsOn5BlJj4Zl2
bz2qDyqSsHvwqbwWAxLToDNln3azkJ9GYg6/TxtaP24i9FdF91lGG2g81Ny22smmBwiUNTUL4jXv
jXh3agsNLWOguqyVHqNIIkPX5/gdLTUl+ecH/HGpXMnQ4zKZuT1ZsVvpIsTRDlfO9P5C7V5/n241
gMu9XZZ9p/KtiqvqHDzUGGQzFl/lgBs+bahYlrEwXm+931gI0p3/yNjQ6zpY0rwmOcxNIKLMFmjy
MQiCO/q1fAw7Np0CrJvRRdTEZFaQ0XOb7KWFh8fjtoQ79oxNmYsQTx4zsLFwissdqyIQERc+sGMO
gmiUgwS07gcRNrVztKOXuejei+BOPfPs/ULBPr+S8XnaP+4E3WXgdzDNKa42g4l8dAtnv1+/BKwk
z37XhT29+MirDkl2t1mMv/+ztjb7LfKW/gbk1TiJA7yLOb5wXj3TilJ0K8VvRnQP11aaS0LJWVVE
sIQAcbfl8inR9YW7x5RwOKPAILs3GeJiSgpoypnpmrqkkRudCkH0Wqj+gR9seW0KEEu/HWnDsLGk
A8tHYv5z8xCGFBq6OWViWlDVbgB8KAznFsXcOuSjWgWakYDmQKl5XyhO7oz1JqoaZ+kc6GbtLnUC
muXsZ93mLCIvVZufL2X79rPMlsBVYISlS0EvMjtA/TLk47wsUWKqyfUPiSLxO8FNcwQoVH+l6TqM
IAKvIL7WF4JxWQJ8cCCb1PgrytjAx0955FfRTycQbfePay4P+bB8B3dHFo8wzIXIjA+7GBNz/lMD
AP7uSfCZw9owLKwhIbrCxax+t+/GAvs5nZMlqlO52dtsYF82Cd+ILJA468dbYBRznyeik3b5tAxA
6q9XANIMp5C+jIg/xzhXu44BXOgfsqBAs8ayuDCjedGPXQJKSAPgFrfKHaI75ey9SpMrdaWfev4p
A0Dihn/AYuBOkhVvWjjOFdA76WDjPlXoCgr9uE6DeG69UaCMIR9YX3O6R9AvTCdRlxNUIto2UXty
20UVkg97n+Bp515Fpkwy2bV1Rfi/MT61tLud7uU0P/yjEosUhX4UuD42rZeNQ4sabfDLproF7Mju
pJ9mhp409kqOHCQm+G/L47uKZYPKH4OhgtzIwG+RjBaA35ewKLKOMtdhK6X0CuUxDlzl+B55X+qT
0ZfzEUeHi+Ngb28AsX6qzQ0wT1esnWFsBw8O0RvBue3+stULaeDFpjgZuCNyxq+827ykYAF2Wc2P
6RpX26mwtRue19Lc3q6oS0H3PwDcuz4lNkUfLbTl1AyP/jhZ5+mf2c6xRIBQMW1D2x02hwigykSX
lLKsKZ36h9Y4s/0OfKajVUWIdq0LoLHB268QERyWL6KkOQ2UE6Qtsr4lQ0MpWAy5B1f400WFJjR6
hufORlUEz4gk+0S22+q55BYRDEBhHS7VfeOXFA6/EXfQK4xQAPvF8o6U9MJIwkTTmnUFYKk0Tup9
IP7KHXjIpGSnO+YmQ2KkTK9fcNliNvqFw+AJ32CbZucBUaBc1VIvCFecc4PwwXiwtqd3wh1i8IeT
ivPLfT1aDomtzgosjQpn1upiZYKt9qwNTnGV+zY/2u5gn5aOrf7e8kl0MUpGwLgaZbkfLKJvpKWU
pTigUfir0/n5ok4tFEWHeUpZcotYBDQtsxTDRMv3ILyMVDWHxRVFYTW+h9sC/5KvyUEVEzfkO49p
JJy++VpIdWpzw8E4zuIlBkyUbL7o56lgOZAnq9auEDetTxvzDlouO8lyj/eltIu7cm30yC4zHDPK
bXhTuJpaWX71BR5+Y4J4xOaqnvVks4UIjRWl5RAFKqewuvWnvVHIc1Lhbz/YSlYJF4GR2IWIwQkH
qNhmA0OvBdNpdjEFKBpdvgC1TU8rsi+uXhz7gXRnEm8i79l+ycdZQDOjVWhh2vLnzIl/STUf5H4d
NVoCfTknnFHhy/s4/xa4K9dhbvXZCP/ni1rYaJOP2UoW6gTNdSkEde9AOKs5MMi9jJwJiJrofjLu
Szawdfh/qgEeJ+lv4+HJYKgJ5oFeKPN3mxamNnoF80b3hlZiwWztSPyaEB/D/f7FuwpJ8a+FL+UL
fqmwpG6Uvm5qxDpRmsQZq1gnvGO0kzxvPY6qKEplV0IbSBPVKCSP9D8Dza9o7oeeIgVAFMOeB0Q3
j4bDqmzSBXc3znWATF7m46BGwo6r++rm9MVzK8JQshaTA627cxJiPIZVpUDzL4OxV/HMdrINMbVw
P+edlOEH6CBLF07jcpZfSYtftJ3YjC7J9MrD1xm/+q6NzxRIx7jaf71PiyBU+UK5YbNRU6r9ndma
n/HjT/D1n9Iriy9KIgtgBjcFuUvrZnl7eutg46FazwYnTF4+5dIWQT5qXO6NFcv9M2abU10hGT4U
A/+E36B3Ed4hgAZurt+6xLZglclkysLwg0FbTGINlOQQXAP5efIxP2SwN50hNhMmUQb4HDb8LNNk
R2xLPsfkTRxDV8o4tMKTjmM6gkXVc+FwAzIn2dfyngBtS605JUv+D0Yam5PmPVGvvrICHUypnB/K
YyHtLBASkF3JH44I5ge4OC4sFVjpfIiHc65MjwbUmSGwd7275SCyHXj4YrIOEG/kCItMUs8ErBUQ
QxbAzFAEjZfnLynph8mTmiRLY59foYktChgd3bZjDJWw/3KwF+yukGdF+Ob5/hJ1xBvIUbLJ+IJ3
nv511R9nFk9HYGqpE0EvZXex2tmoWcX40ji0t/gCTpf//qUnUuvIK0mPYJEM3kBEbasRewmJTRNr
wk5pnou+o7EyIvaa8Vd6fz+wvYBuJO2TdvJTNkY+Y2dTXuUMXf6EP1HLmOqiIbgwDswFisQqCDCV
+wTk2mQ5OLzYzPQL1jJ0k/D4rLft81g7k/n4eMm9zraPH4pWKEmAw+WQxKiizDjQCZtEYfh3Ns0o
+q6Hu/IOc4X27G/upCdr51i5R5+k0AJygZwQWp1ssE2QLqEiizn4+/nTpxQHSKmvh/AEQWnqb7vq
NSY54vT/5AqOiyzfhhbStk3hrO+Es+K/alrgTS5vHfypeGt6SqSEtnWQVB6hRwud6BAsSOE2mFJK
r7WDOAPMeG/v6vL36Ahuo9k/eU/ZeFFpHDR/jdMSxBxguFy6fHuhMcM2A8f2hT7gpHhvhoFdl/d6
WxVLEvULAklGc3Q1NrjLGpuXGrPiI78tqjXSfpagW0WuSVIX8ds1mCpDuYrDnhD5b/A/0X4ZlBDd
5XmXxn3v2bTqs9uYYDh1zaJ4EqGwoTb7XZ1va4KGQ5kDQ2KO7qGjlglo0F2nOggYXrmUdUHYR/Ac
aj1X6ZctpzZiNa4UKeHY734UTHPTaO0zC0ueOw+EXWVsu7w5QeA7617EDo3du1u19SzWRlImgDtg
qASRnrBys49FAnva9fAsOldaeQOWZ76ja/7Vhgjz4fqaHdj7QKy6u4kTu3zG+eqsKHFIT1CBjW+A
xFqkHKHOKZ0J3iWepNCAPP+CJmYnjxyPYf/cgTzsK4nErTwj4Lh1OhFdW/iqsNcqEhYMJSvbX+W8
kMmQ4TRlUG3iBy+2RSEMpeZxvJgSfReyMLJjogwZm79kZ8ziF+8J9GzqebT7m6g7YI9jEg/v9dHM
U3pz5MDZ9xaCw4SM8bHwyPQPXqARKxnsOVC4RcbY6HrxJ4G9ZCvf7blGzk+ypmSDlTLhY38BmSRr
Qa1Vxl8mk2R+j25r4uG9h+veH1e0THfkzybmhHEGlaeK3FndtdDmv1gII600L5toIycPyC/2GKFW
86rQqZG+EbccJX8URCyVzyall/MMpjOPjA+POJoZPqK4AEPkJbrYlcO7yonBTAHchA+TtvRgBKph
yaTOFJ+NV5jiWiiLgeNVZg2XYDExnHYz87OzY9PZJBazD8q+fTc/7xLzR1LPFmBvmTJ8pNsxTg0j
tdH3HYFSW7tjEj47gCIvk0ZQ7UlLzi5Wv8R3oIFdeC32uTJ+diEZxjXtIBIgiOdqLmQsA6R8OLQ+
XMx4ulMC0heOnwvDGt5bL8HL2SpDdTsk+30SJ00adsPHUzLZuykYThaXX2GB1wQaGepJiYkiwIwW
pCAVfB9/OrPBR9fDrTHH0qbVaEv/jz/0oj9VMDW4M4qgFXJ0oiXsqGv/k3zNwBkOdui6IEIsmvtZ
n3eesoyhqWLpaWNVUFpQs/mKhmuOQQrhH1wREsFzZo8HMaJ2WOhc6ig2vWjgWpAKMaMcbj/UBR64
KmXhmmi4yjDxC/M6aL0Wr6BE/a2tFNQhdVmx+P2SoVVHfqoWVvcFfDbGeriZjpViJvoAWe837bSI
vgE94qY6+zgfjIV/4IEkQnm3D0xpXkjM+iZnQ6DZsiBd5hpCuUwpFFxd9s+YAhWCK6pRQFuFimru
4XmkKQQ6cqSBZ6i0L+WMup8e8MO/5ZX4KkgjuJyXqJRP1iRaeocNmtOoWNO9wdtKKFVLo068fbFl
8h/Pfeex23UpSUCexvX1CX2YVXmJ6e1lh4L0/2CUfqGBFqUFrSpIQDoUjcounC8SWGWcYPqVOs3Y
F6xqV/snY1+EHR4wVdrj4asxN+WX+F4clZHLHnezYNz+5UWUc1e0POkk3BxFjjmMi8LzXfHEapGQ
tOyDPJN96FMwEwWmqubQyhblMp/kCxmEMXg9tziyOYlpHVl6hDpvthXB8ugc//KOrrdu/DfBCTlI
FOH3eNlS94r2JS6UK4rFRLHjkL85jNQvlDyr2GP3NTSBe65dLmjUrBChhrIbKGKR+YCuwzVatsBU
7bcPVfbXCvqabvvsKJ3B+2Avzdrh4TL9ukfKLGiNmXVKrvwz7t0JPgYrUAbhSjT2QsISNS5ksnwq
egoCdUq3MOltl8Onp6IZT5EsNGnc6tav7f9qPWwVaYHtZwwb3F1xIDSC+bTrHjKcdHeooBTDgZZD
++5zKRzVpYa0m+TBoBmbx++o2p9LRB9q5TguWDs77GRIhdf2AGHNxRVjPgvMnQ5LpE/xKjyxmsOY
E6zW7yQa3f87PHRJ8QFa+itnA9rdxUtXXTXp86xX3r8RY+V7tWYKaH4fRZ+FrAby1tYk1dPP5YUu
tu3P8TL1jNDPce2RsY8xD+2CQLpS0UT932TPdLfouuThv2LBf60SjGLMPKDCsLbfenn/whagD86O
Y+Du6HuAoSD7kDyghwCgpq2fE6HsgC216VUYn+okxbyndEzLsOj6EYgI2CyQHehrcUvb8CiC4TSG
+cYcjLzthgSbEZPmcfTcmps3YiwkKRBSYYBvNlSaaVrV7zlSrJf6LoF2PuGwOIxVDmDMiRdGWExs
YtQRsZYONppEvvF3BQGhOmRJIrVPRnTto9X8j3sMrk/4kVSjlWrbVupanPWLJnCBmEKaCQXCSZmz
NM22j/B6I1JDg1oK7BjyTAnYo9/3BFrwMQTPfwfPrvplMVg5DVwkUOHhQn1h1uMKFko9QzJ/eZo6
GTO5z5IU+9ZskV3HJssBcUzCwxUc0U9tP5rj/GN0gc1jzN9DoIixXpVJ3iy0XCOSnm+ZuxUkYfx2
eFZLLCSsB2wEaoiHRvs+47gqciXtKToO1eTWak4rECoK9TbLSGSGH04/7X2Vm7Q+mp0F9NpaJSJU
Y7GqmbwP9EirY940hrEiCI5bsXDSKibynoiOzRlrkzonBEAFKrEo4vB2e3COkLkSs9WiQ2z6/lZv
yjhzFmZLKIRJ0cYtVrFQnZH/0FSl6X8n0l3Zhi5QFLk6Lz/8Izk8VW12gI4yLeyG4tiAKF41dXxm
WpnbmBFzRLsrpZQMZpifkBhdT9Ets4w4khE4vpfMgPYDb6DK3y459bFMVFyJLUX7xQILXC4UGjYm
79AZ8pu+uCLHVuXIRqY0QzyFYnw3JCt0/bgEuGophHxoXNJmXe5sjwcFcUSjDZC8T27okQdOcttZ
aypeoLA+1L7w+jDjX8s0qC4MaCjxWLv3z3agMwqVwEFQbMAyycyUt/fCMIKdts5t/LsP0g9ZMK1V
YTrGjdogA0PduxifUhlS9IPnAXPpeQ6uk9V/7bNWdMp+yg7l86h78F5ILGYrHHi8UD5B7AHxx6Yv
Lbdpt9uNebqadNlSLyOYueATuY59EsoPKNir3X9e6TdeJrBq5DzZak23LDFBbiVPseOAlGZFwoAB
zmBcKmyQ63whoDn9dKpe1W9yYFh0booMwwDrbjj/w60EWFlNMfP//1w+L2Jw3ePgG7HzlpMu0v2q
REqPHc9zd7eVeCJZOiss8K03/TZxSZ20hIfjF3D4x+IxjiyGEQi2wTmAh/IWyFVxmxyhjuxPm/w8
0TC3sBiJlHiiTNQfzfsKKe98oTuTg6ZumAIpoZZ1GpxRkDhupLp5rBcmQLVjYvXCIyDTxLM11VcN
6zZ4kqMRfXBycx/YsHVeFlB+db1iYCVqlitvkXUW/NgHLdOX8gwznKfEcVNfCpDljyQqkK+l3oiJ
dsijVIQYmyCBXZAKfN7DRANzW5eDlOQo8ywbtwQaDDh49uSLPFP3/a4ORJl5za9oBxWrUbl817mP
SmLx4xI0xJMSLKLVJLJ6ebTxlxQ2gI5hc6oIlkqxPISeLljHR9Q17XbN/eHfkqVbL4lPDfiu7kis
PPFZE0JtM+P2Zd47SJnkr8Hr9xoV77yWesQQW7t9YD8DnES13CmvVTo0bMU5TJ8ZbAXzdiAaFH7U
9XHAG2L06guxVZ4SMY1lIhlMj8/ryFrYW30VqaBt9GNofMsjHaayozpKW+KRXie+y9gve4tRgZil
KZQjNNFMGizqDK7nYp5/9G4kabgrxEkOzo7mTJRZ5FOQvIhWmihJXiofD8Kj51dfg2MIoOTWmV8J
yXXsrxYUs/yXsUHaB5bY0X6UUZTTKycP0wgM1AL5uL2gJLzJh9sck8/QiEPRk/SEJQeWi4egNz/P
JVlJ8pikHKGC/1zstgkqDep8xAWmfPBzNi3pW2Mt5JI+7XyJULuUdYXyswJ6uZX38Xe/tOlfnjQH
w0c0ceQMdr0w1pG05etQGQQOEme7bXdtBEoyjFnxXSuahLqmAUiGPm18Dq2ILFGoHduWd5bdcMM/
RDwXJ7VOifRBXl6JrWdgwObc341gNU08ciGo6eTnF0DyMSVFVvuzdDo5owSiEhU9fQVVNY9VFTPb
yhBDJDrMtNeIh5Yy+eSa5K6BCWqTnySR/iiksBDIo+21HGc7Y7lZBuuBZC8AeyV5JfMqxLK09WcF
0uxZljhKUPkkMaoN0qckvmFNPgqykP3NDEZaDgmSAL5PAPgOP7upkylSCRJS5jRU58OVPSuH9hsH
zVkTUvxEEtNO1A2ialuim5w5BgmqRm07Ucbcd9xuteJdpfagyNb3BLBcPWAuB5zy+kJeMP0O9zNe
dE8ectiOyUKtn03j7/Tv4Q4o5kNHPnzL1vWWh55TA6OvB8dF/eB0rADxdgzydS+6lH+n6yGQrLR3
gS5sVvUz0918xQONtQkdRynEY7kH20v3Nh2C3Bkok4z8HFOa9si3AWnLyArryB1aZN3MgDMdYK0Q
pe+dbbONLqICU5Nx8kSaGRxHKlwB0rE4gwLXLqLH9b/K4PybhYDQ7lpgCc4VNgmHbG9529LShLVG
ZVCavoJZH436WDGHD5Q3y1XOKixHyHom5EyKzY+L9vIzy+ju/mWdufnQXUNjeI87HRw9gz8m32p4
AhICimR2YZjfKYVeACI2OubZ2tz++Xp63fP2FpKLUhrAzddL3p4hnz4KPbuB2PiHNnkorgrqghRR
2TntOUXcdn548AN4YrC4NubJiG3pxYqYDtRlh00iD2Ni6lwJwv0vjSR5nC3NbMMaHAmVoL++O+l5
k88uODzUeQLu48MD9UAe/YBFZYei9GR22+wqzImSZiwF2mHtTf9V91PzGiBhPpoVtL2jMJZk4ccU
rb/vu+p69AUfVoL0KfXvxqb91GxaDetOIu58Gbw+/Dpwb/Y11sc63Ev8Nu6QjNagy+QwD749FgEI
nMRAfAkUlSH8Osmlue3NRK6zgwO9r0/bcCVP0OhpIMiZ3PD0SyqthV5W07Q348fRw9c+ICr2t3QB
dVf1YxKXVJo8svbFThwqNSJr13jHHMXbyY3BpEcTuEzgXrE+63UBN/f64SfGjGUio7oormas8lvZ
S7ffgNq9Ju7XHKL1NjRwjyIueC6DQXZ34Qsj6RFHKNlUE9i9ofE1myIaIuqz1NUYDolKUCNZQQPD
uhFyhyG0vY9e97IfeiMIHDqK+N/4RqgoWuAwH/yF2NDE2XKH/YBaLHD+RlEdMMaXbzA+//vHNjTh
AytEl9rmfiOWxEA0twvVaiMp08CzzwF6BO/Y4z2ZukQpmfoclv+/CFPtFVT0GA/1xlmBa3qb5Kvh
8g1a8oWAMbb0r9rBFH8tpmd0eQqn5QcfmA+djCEehjVVsC50QFO0sNwEJ9JxAjMrHnLuSBbj/rLw
s/U9psY3gWxC4vnTmV6dL86p9ZHAMUZghyKy69ryUKqK2udoo/Upa2xzXNDCY5cU4ZxxYf7X1PPW
akgacj9YsThTwrg8rnoLjdhR9MC9na3afcSfLbS+OGjRr7wlg1HyOYNI5Upe6AM5fq8OosynWpNi
dtehmSnr+Hosq/CKyVTX04JvP/xeoSh5fqpKxgKi20LGXFuFEosyVR4ToaGl7mk1nTq+yM2IhNE8
l8LIDyarNGmfgSwDXegL1f5UcJTmaIKclFOVTGyC4eQU8fpcBEuSPoGZDynm1N1qn57gNHCOVais
uEK3qwXWERG/XVtva+Tta/o+ZSWD0Hzyw9FaygUlVTHUFpmc1EgAMuxn8uM2yB/MYct1cawSUw2j
/7LHqUrBf9s8J1JHU0ifEc2d2Tq2SKqmFvlAHb6ojnJX1tXQkJrI/G9LubcksGP9zj97aHk39O3R
4a8pcA/Ey4O8WytTWFVyyqaAwwdnp3uIrVGxqp36uaQKp1NoJ5w3qNSjHSZTRIjcv1VtBRgnO+pN
gbG5SlD/hxoqBLmW9Efz3HFp0zAKr7bXBah198SeExiIhsIRcCssi30Xb0FnL2xByCukdPE76+7a
v2YELkB4d8YmAzdARr9gi3LgPSFatWzV1wkmfDZjWiseQBR9jAnp40BFUuHAO2pRzGgA3GgM+s/F
rDqgYQ8wmzC/ZYo1MvWPMmImJZiItMKY6QsKGaAXSrCASxLVlN7achemw4CFpX1ddKN+E4dZt4Pt
X/qQGN/VPzGC1Cbu7iAEMi/bYErSzg8C/j0gRSrnmC8ItMfgRAAV07L4CYknTdf51oO57NvKYBWv
e7PWozdxKbdC1utjGa7/XTplN4O1glec0aKaxA9D6s9lCngKlSfjZxx64yN0zQh4BJ7QChShWvkn
7eB+xLFHHAht+dbPfsCAqOtcCN9LwakVa/NQPpivj32kYHU1/beLYIl0/3NgYSO7kj4AR4+BHzwZ
E6roeJvc3V7umEXoAEd36NYUUTki08LHQ80hm3FAxiFcNHizpSxZP59j6IeaJNdArbVGcT7cU2np
nt7yfApoQ5r4pfkXL/CRqkt7YVnzIA85qUlmcfzvPgvJR4NysQBarQ9cdy52z4ko4FaBZDBX8ejB
MnKreS1zpXlkmMAfQJ0J2R04xWofyPKbrxw0kMlMjw9rSee4lbtq7Sizof3ksp46S8I6a1fqG8Wm
DP8BpUQ/KrZfTWNKdC4T38KWmkJmbP6pamrK0kSL8jRFoGOLaaXYolqlaZ5OA0sE9sytcM+I66Ra
CbMoKBa4RBE1rXHDMSBvkbQ2EaCYgs6EKE8XvYESxKBcn1pN0d9a1oui3+SZIdSc7stylF5+1O3l
pPSjXqw667YDg9g6/oQ5PRHUmoYWj1Lh1rRE3dJvv8cyN+fK3FDZXCr7HfSWSOfW1r6j8yZp9iAL
DEi2HJAS31VFQzHJSpMdrIhDfELQltfHKu1N7oJlaOFk//USfi92UKsdQ0K5YiQ2/rN2LG1fTPnj
IPKMDodtVmjITtrvsXyzPlanXqDV8An7YDhCGTT4OOtbpTFwguWg0pMrrSbwP7XhG9n+If/qMi+3
yu6ge0AaBQBevQeBf+w1lzzoVHWBgHShN4LO+pqws5h/Y5uzuIPbDmxVp5z1hm9dU7/EE4SDWbXi
BIHWgJ5T5saZrAI93J6AxcmA2jlrmUuMfMfRKw1GklhxESQKWE3hkHvyxn+pfka796QDx+Y4dICx
QDILot16RUeZlOzU11m7FrnREMG0wQNluyrr04h4LNcvM4ZRooxKwnoTt9W3CxhF9Kxbe7E4k25v
W2bh6aS2PH2scxeDwUN9IvrAJnAe3RElxFfhiOdKsruXsz3MNF9M2TuxpTYWfiOazyjA1mcQtLdv
GwL5MKsMPLR6mzg3klZE+T/CNK0D+H5ieTAe5vKC+jcuNcucnWnge+X8zFhc1XnlTNuWt63qYSWz
WkSkquBhVRnH+D9szKVqFAXlW1WcE+fBeBDHnRe9agWdfKWvsfCe0bPkKdH1Ke9LdY4zJ6UVWiA3
YM8fIShI6iMx0frdp/JL+pOf7mSzbal4j0nYqDioX6QoUyLkOhAnHrjlmzvT+fB9Bg76gOWg5Ecf
u9gcko1M/fSLupE5TYERvitwfaPccfjABcDv4v6mhynM24F3x4Qj5JldURIonRuzDkvzwtaxl7O2
/el2iP4lc8AZ+9EHnRZuaFwaYQTx80eoxDLpyXrIkaGj0rRgbtqzPabQ3YVQu1gFpxhSprZVfC72
Ee9lAenb3AyTTnPXwHCT5/YqxFclEphK09zFIjWoTKD2fZ0kASGXXlzql8q0YwjmqNY38iOTHLal
/mM/9ErnlyDO31bFESh6riCC2xXvlODD6qMgaJox03mTe+/UxOFr+Aig924Y3vnnsVBI/c4Rc58p
BDDmhaKFREGwHMwxOWoCdn6xctmcCY/eJ0kAOtdW3AK3g0lv3j27JiR0zRF5f0ZQ8I6qrkNkH4ow
H7xuhTG3xT7XFlQmPJTzEiv7rhfk1MHeJwxXugBCHWlqXVv5R+z0GXJQw/eEBlGCPHB7mD16J6Nt
BIk1yTBMxlShMdW0GrHB72rpg21gYPGCy5WKYtzFg5QpiJP5TRguiXiegMtNtPR9M+8QMoYAHtrd
jK4w+eXlfe34uFlPeLnPxK84r6M8wkL3e+7QnehIqAtRPdV1y1hPz2ddhxgp223+D8VZ6c0fm51z
F4rYSZQzZjt4Yb3CpjRpb10GHyJ4SK5VRtJehHJxu3EF44Bfm3cHKrYPCf4BFS3z+YamhGEdNdO3
Tr2wHiIo6J3XivDgh5FqcnvUBAmbw4vDSaQo/EFsvuHlNaX9gLM35zeX202A6DG9JyDjDkywwZZG
Al+Fl0L1ykuQkVftizwn01rG1N5jzoMruEsc/tlO2Yr++Oga+pvWtnsaFnFdlXYmPtrfRjhGzLYp
OHDj4tiF46CzTWUfKZJhaGDbJ8NQOdrtgBgM0WAb5cjojP9sp7uhdLtoQfS6u2nSHdVYTxbcKMHP
mj0f45+QbE8+Gdj9OkKjCI/kgFQylXD3HWp613Zj8MGyHD92wBTbSS0xkDGwsXYd3oHceRkHj4Os
D1X9ho86hFdqBx31D1ePOdT1nSJzbgkSKFccxoon41zrY8fnwMpMmexTnxRKQq9zKdmlsxLtbi47
6NyrRXaQvg9VArPnOpvu3dCr43VgUjm2cS+G7ZOSPv7OzoMm/6i5imx4ZOUOy2NOFRwJWAhSVzoT
5znLQHybHClNpbxlRI3hw6Dyu/V9kO8bxRd+vxrG0ENzW3jiaD1MqlvERVb8Vn/y3hx4Xbrql+V7
AS/gfPy4WwrmR1P9Cj6/JcHQeRqlnQTAVpL+5T8DMPrB4lhXYNpZ/uUmdpAswNojo/YTfAjnx9em
RwF7+/Et9wjRdWnE9BzD3wXJcfKWkfIKV9BGOcY0BVVgEw6VXU55kpYBwed4ufs82gwmGuNud/Rm
aKBGbQndcUIcXOZllXMLe6wpJ8Ja4rEEHBfHboLSDugiYQKBiMj+JhiEYfkrW6sjokcIw6XP3cBc
jQTfXrheg7AcUVCeEMAsfnq/7DcgESWfdhoh+3D+rlWOFSWpSy11nK11vIK6vJV1c48fXwOrpai2
2Wv5FVvFueQbm+Bax/iHQcWNh/8WTZq7wlu2ruFWEbywbSgqDWPdIAI5ZuuCEG4J9cZEr7C1W4LK
UurwqifHB8jfAFeEQl4etWIlQb4ucPIW8zmVpzZ3H4Ejs6J0yM7S27OIqmJUkhprNg6fo8rHJY6V
rzp7kW2h/g/S4Jsw3FHGgCNUbI4VIAXjDUItOufLVQ/6MU7XhlwKsiHkyT0Vz7J4/P0h7oHoFych
sYycmh9Sx5YdqNPUm5o/Osi3W+SN0J+Y2hV6UXhAtXaNm+JseP6hP+Avyg9NcdF2/L/JXUP7h4tB
EMlcN0ObJqiL0AE/OrM+a4to6wif1z29b04Tniw2YqwhhVbQFrWGE1uUA01e+8JvKe2tRgcQNYPf
qD4OIxbY6apofWhuvN+ciRFVuXe9HGicRd0PfoN1QN+VtWmLEICoFaVT+mYZH5ZnVMH6Q52pRk6J
exe1s4EBUOqFxEvWu0XWONbz4pwed6rD3RTveEKY+bjICRXgZiniUOzbgBmXrN45JsFKK9UKxycK
Pa7VP9ce80fFpvZPho/r+9al3oOTz8UtN47lkssNdpvJJdNDjKzHVOe3UYfd4cLCm4KmhWBtS1pL
JXZMzURd+Ssd/3psmYJOEFH6IHLUkdv8MZewU4acfX+mPHgVBMfjHcuZtdnC/FRkR8qe6VpNFLsW
m40z3jBtDiVaABNiutO3XM+idHCyXpqrbpaxhezFwqpNJaEVz0w6SZLV59869bs/LBMLaIU6MNEA
RW1zJee0WxT5QhrQE3rXNEt+hFqXU6kGOxv5dHeTRoN1QDwCpbVl1VGVdGiUdOLeZ4nnO0koSnt6
wC5bMzBU/fJwAAHg298qA0S1iMuH7LhUNNhf40BeEKTR2GyhfqIFJ5SVPBPuK6+P0O6lf3G5yqQW
1IMDbUdUzR6xJM5tW/nUywVdtBtDgxoB9X3dUZjnCv0pvtsxTzpEO8bAX7aU6Gk6zd5IZGXMU6mx
i5Zrry4v87U8tq1JV2GlMO/PdNG6zWFWBkuzBI3jWQwdGZWkv3Cuupd4OpGe6fBNayh4P9nx/8W0
ewcJjv9044dNYurO7kDaXp002+/pY7CNXNQA6+dAGo8/X8Tbzrqw3+DQIF4SShCSjKO/PLTTrDrq
tQvPh79ieRUKw2wUSTriYlBkHeWz3jTC3R4QQYOlAykvGLF4An4Ean8Itw/MQCX9TnUzS5aKDnJH
BNQhm449CXZ+KAS8xruo/NIvFs5k7d+xMzbpguuSHfsICim59a7VxeOmCaycOQLdLCdDCXAk//PP
UiqcGylsWnigerYIX85brGNXdJ3wd7gxx+iNKh9sggc7v+tPcWt67Qv0xVOAnL7Jc3ezX6i36+84
z9lKx8IGLgxgMdKX4Aw6MWdIxZgL0wZeWK3KiG8SBomlrI9Z1600nBpWYAIhKib7RvYOGlX9JNDJ
L6dSR4fSmED1ReQH4910kMFAddsHKWux/RTEKmvJ1NDmMwAwA7kB+ZcsuNN920cQI0EMI1Qk3KB2
zY6E+WWiKEJ8aqqVGEzuflEp64PXIB7gpGRDDLcWqZShyiNXPiISwn4+8YxLntuqR+0T1j11UcPD
vAAzssVPbpfujk1ktFS+Hma1A8I+KbbJ1qfy4dH/5WnYlY8lwRVlkjTOyY6Z2wuCEtZLqFf7SO+z
jbGgDn6fNekm7uzLHoB+D52/PGwYLOiZkRFcWCYQGWEtgDrpoJ5bQGDLWjmSXnQFGJwDVIwkeojV
0kRzBRR/GNdqbCjiPr332hVbBrHsiLTnwskl80IWjLlAx1s2AV1e5pT8FV8PgjhzQ4wxpJ6M4515
m39CHhwv8pJoKI7C0+ZnGiM/tQI0aL6/e3a8VtiU/4aNgCwcrefdKEkWLZWOk4Lk5zKHKTGoYKyH
my3kTGls5cUYbJK/kGXT3Y+qzrpXacuRp8m7Lv8HsMp+fcm7CeKtEPB4stPn87m9uqROBWVGyuT4
kpWCtT+fGS4Ir7CAkFgM0EP0bkoFjh/yCBPTMK/TLGaFNlpWPKywn5jeIxr/3tOgyRZnh+oyhNYn
rtaeHklGEsnT4ppR0/LQoDDA8P+ccv4wBihA3sGdIbmd3hQN/ohRSxPBkj3eyzSESbHNapD3b94q
e0qMGcTIflvtAJh6B/tbvDZBHJ0rL4d/kFzsOc0riGPHKe4pn1JXN7Q6kFSt5hOxWzLwPkZ2sGEy
tJIe+o4CNUMOUR7VMG8Z/emLb5JrhbRfqvtrtkaO0VLHrFyZwUD/5QeTwiRj9vcm+jaTuYFssEIL
zximDyhjJ3YNR8b2vfTvvI+N+xyBsiMXk1JEzIqgxHu+X0IJnn8Sfcxapd1ElDP7EWkpRerg8rze
J9SYbfUoI8+BuKBe5eD9YZ4yB9+UP7YaDsa/Pi+FTp4KHxZtfQrtOpZ9OBF4Pp2uA24lIJKcWGit
6EaE7rEycvck0sHF5iYGhD40IpNFcfiSKLgLKd28C2Jr94n0NuNzorqFuOQCCocahtgUA7UFrWS2
/RjkY1FhB8zmTGXgKbJpfngl26c9QZVTsKK4j9ufxIK4ujqwpxGG+UjQi0ssprqJw608djwi7hzH
TitlEn0D0XAMuLt3Go0p4TwmmU3Bydy5MgJqRtT1cGYnSvpy0RUdlU4lN6M/Hy3G9ViuZdqp55DY
VQh+CjpaESLei0DOLuRamQNID6R2ZuATnGu5GjCBkqCbdSKNMumzV9r5SwcNt8oVXpaHj222pYta
2e+PSb5FaOFesTrFaIY7eO3tqJOLCTq1UB8vq5SkDdqZBV6InRHvH5EYvM0e71un8ag93zIyxCfO
ThIHnP04ifj/min8yAsoGX2yrGxO+zr6C0jePq4D4eNXSGjqbKJd2SUYHSDmazEltAsID94JXFlg
+jyOIgMZMTzQb5LI5KHw0HuOKk92BrQbo8bmvbZZV2dY6h8ikeTQlXbfPgBKDqL4NsG2lAGpDXTO
6xSMHVBHXZHg1oZrxDNxuP20DHicB4ZbFMHV77NXPBF+Z/w4QREm1HFNpSpip42MkOHP9y7k74eZ
gLROfxeBDLG86X9OVOfSAlAk2jji+oOcbqtpxQK7WfOQgi4WpHzRyjjduKNCC8ocxiuTpY0bgrUb
JVVqxH2l4kU8N8uHoW0VM80ZHvpQfbyhXc3s3+sg6mJaxhbr+sjAszOWfT8prjRR1i96xXuAlFMI
3P/aG7sWZdVnYE11vO5xJs0nXAU7+5wprtfMnZO5vgz16+Kgj637xHiZGPs9hMaj6SvTcjdq0sv5
C0gQLzUhMcuW/JItzoSCumZztU5aMZXRSro5CIF3fUsFaZfSo6CvPXHjFHrPo0ShnjjI69uvaAsJ
at54tsZRnqdPa0NwU7u6oa27N1DP+RwbLX2ts5rI5f4Sq6dQizFtviWcRWGZtNfEPYe6mamcep8J
sJFpiE/K/jZNv3cfl/QRMgiHn/Y5SE0hfxBfNOszsa0lLKA9eazb8vLTv5kM8Wmr/O5pFnnwFrPq
A0JNYNtDjpb9Ynr9c7yLxaeMGTumfPAONJgE/4xiq5N7hfEBwU+3a8Syh0mBOKJVcjKyxNKAsH2B
ZW73bRSUgFQyacucUXP2jvxtON5YDJdVHqQPd88R2h9Fa0W+Okvi0Sqyuh6FWEQHiIusUei3o7Rs
6PxXdsmsNSMplyTwrToaNa6iRNI9TPeUvCMHbqRjIY2KngjIyQRPW3UsiCZIdLXuEnxlBPvhuo12
s6Ie3WVyU3l+swsKRAkZQc3o9gmdwbWTRBJii9vNJr6nPNf/k/Lr+VoVr03XBGLHTs06nFREgrKP
WsD22zUODpPgcBMiS+Bf37P1CIfq4qwzmJyxMOqIHOItprtslGhajOjvq/PEZW8G+XZf/RLT5elD
W9pEegwnHCV66s0rRRYz9MpcR9iwQu4dYu1vAhJR/+N23W5HdeQ7UGF42nMx8T9OsiFGRSCLuafA
cjZDj2vJopkShezn+VR1EZi8iMKYPL2x4ZMBBZ42hON41GvNrUaqqG5uKTgSLMgxLwyEfX0JqAKA
xAsXs9n+Nb+0bnMk7YA50PtMb6tPEcy7duZoyN+a7QAotbykGm63D5qI3MWfnPMv7j39RWdSA+wz
k86fPfZ7NhvTsFjBrs8iPCitkaLopUpsRnAFQNS3bDlrQnvKlZo7Edn+Iy3XVUdtofzJnk62110N
JTMdoctr9HH7kmTxlQ/L0rX3m7v8f+VOUPCwhEoo5wMlHbjytyKQDhUlJkCwY1uGP86pHbZMU7KL
ulE+qbJtue+0qLgo2iZLKbFit4QqqQ+0MxSur3HLGPWwxGkB3xz1mYiZSYbFADuHbo9/zHuL623M
3C1xeoDTmZWq/YvggdHbwmfPsKfWTsP9HkvShO8A998fixI5w2V+3/BIYou3JF/leJSoEJ2zev7W
scFwUXm1+4KX4skafzZY6iUPGhbdbIal71iCOq3ywd9QDNQs0MIZ0pcDC7hxugaWCTo5GKyMDenJ
D2J1mZOGhCfan6PR1Ccdk2lG10d8icxx6NgaI2+yeC/ktHZxyJEn3R5zC0EnZq3ynG0f6BU8nIHN
QZ3oEJDdAAewwNqW7WKAvEZWde6mxtwLpDn41tFkXy7JX2I1PsTlXD4KAwImGMt6fo8wBrxjopsO
c8drKQbAYk3P9KYqB06bqG+G97zTzxYbCoxvCc0m37Nb+RXTt1iGmK8G7MoPj7o/ojrtl3fUc+2G
IjXeJwB7Fs4/VnXskTlMKUjywX7MI56gH4bN49FZut1rj1YJsQZ9Me/lTo6fWtkjeff4m4uXM4ma
OpKSozVMIprzjPkvm+FbL0RXOZ9F6DryYW+lGYO71fzk1eHJGyzfZmKQ5sqXSUXniQEjCPMue0KI
58f6F7QB8Ymy+j7wE3F5JZT3uknrmlBlbOyz8LnVOJ1dUKsrFyriJE2yCf407jMIanvc9TWse762
Agi8bknPqzSdJvX7aIRuh01lvw0QmxA2rbJiGXoNpr6kX3WSqo51cjbaLXW0J6+wRMkdgEzHPU1G
Jomfdrfq5oyzdqWtnDsRHJ0zMHBP8Ve+izSt2+fcVZZtP2EbhPxCYd9SvNS1LAEJ7Ww/tcp21MIa
fqXtWANSut5SX/aSAEBnNNfH73sCeXduHdgYJfzB2fZI0rYMWkzwdsLAp17V5dSyzRPrbmQKM8Gc
7UvShppRn9ELxgNQdbe4Kt09FEFjj7UbA9ZxkyOkSj0/bgAevTHEzV3AXIAvZ7dApCEEUGkBkBOR
MdpzTNqJbAEA7bW6C5leb1TTKVpOmqMSaC5Kg7EjxZthPhzPL3b+qBZMyPlhJcK9fB6gX42+oNG7
ZUIOa8Hfy/fezppRagthcT07RoXR14Qmak9NHuACqMEUiYggE5AU2jzwxf6A43ZJqtpz95NXruRF
XjMacONjdNjP8LX3+RAI5pIue0F0N+/r9eZfkikHHNkUkMA84SVsKweObbijv5Zqw+BD7k6603dU
EwLFfBdSjUOAIsMwhyv0vwkR4+sxavU8CKIa5lvT+NpQusRUKrSkJv235yn9/NheTRq5256Zt9E6
6nK7nzNHWPEu1DUsDnQ3cS1WIRzo+KvoJsgnSACVLEZDNdpqc4+nkc4g/qLHS1Ri7M3EsBF4U/pU
cu9ngKzHSSrJBBkylX8Km8Xv5UtIeT/6YZyrOKMBa8taJp+szReWZKLZbwSE/V5Sidx6WuLbXx0e
vWUSjXBWneUWWzrI6ybXagcahhSuFQ+KVQUPTEC/dhbLmaRQuKx3g1+n1Aya1JTahBFTFInwgQvh
kzxAASFrzbovOY6ghpudZIXAzI70vzK6c4uvAJR6u1WYLQriOaPrwp4FJA0y/EaHzVafonZQCPiJ
t3hJTSmxqYcfG8QDdjbQQuexpzo0mzmVrCkyetVzF8kHeB3BWI/DhB6E3n/FUIy9+72P33POxBkE
EcuPOMeVes76JRGOsosXXJNzYaIozejhslckYHmIxjGcRCcvkzTUT5jZ1qgffwpWpbVnq9GiTBAg
801k+uUxlLtFItdfWIN8A7rNXXMoIKw2dabGtvc90Bep89NuEBJRuR3tR605G3Fd8BpSigKu4/5b
ofixRcXh4gy9PBFdQdeYUIIDJszMr92zyg9X3Mr1aLgGRw2CCZJUFi/QqzJ0whGuCbqIJaczezkP
au33NUcBCDvCQGB/U9gdiovNIXR6AW7ZGaVlL+40AFqHgwFuQZXmcjGA3sbOv1Hi2rMVfb4vNhbj
C2nK3ERgW6SzyPancUv0KOpzUws2L3wCy5Jlkv7jpLbGHuJljxEKRcFMgPB8Gk/HLbrBmpOpBDzd
BkNuMnfI2IEB3cUC3wqDjfTNygkidpet2GaMCjKi3jSZtB2kfjS1PjD2Qi8VCSFAx+k3IikeuX53
jmYnIIh6AvE7OTC3HQtAshXAMonOqOoTbEZzjBA9CRyE12LZ4/nhepHEkbQrO5ggDkZj76ulMifl
QBOIf0BmZpUZYZfVeWOpIl5co8LdtG/vtFMoXOuWzIe6ylLNenWOAyiVYP5j995eNkLdjqcQCfXB
u3hWG9yC2J6D2x7GYVjyZI3bJ1qnxIeRM8uVgFsDbQ+OoQRS4TK+iseM5vokVTn1GZW9W+1+dpRr
L1s5oawGD8lKu5T2BJl38CLGBRWLZSr/ApRFAjfhwI2WfmXKHdfWcz2Y3ewu25pZfOQ7D7rC0NCe
ngJiAW7KVA7xHDxSCrRPIsR7Mv9l4eoMNuKk9KROFJNNa8p2iXRa1Vy7DNsWfskOW2sTG+KlsgyY
EFXCb4imNOeIGLuQTb3cdUfSP0knyHYu9WjXe1UC35/JtnUUorSo8zmIfEU+QyjZK7pbedXo67nN
iTzzsVEbl6mEPBhValj+2hIr1sewMTbLv7jzXXcAHmuWq6XbjEZ35sPUc87LLca1Aj+Kbet/BWh1
SxF6HeK+Mi/VrdiCpMOSyo0lKzYMooPSCwDcfDgvGda5DGibf7G2ssHEl+kwRw4UB/Och8kyC5X3
csOHMa6ZjRCF7VvDqXDUnzsJDqtbcFWSrMFkCdrQDSV7E+ONYrCIYodFT86elYm6TRpxipA5mG1E
TzZsp3n1iDA1+FcNZ98dvxpg1Xd6TJRnTSwQJP0yhZIuu9dONjsCfoxmI6E8+RPqV7OWroTkoLZH
bMP28Wp0iAjZ0M/mVu2eibUeTYDw1+K+Dlc/4P2bJwjCHXfXx+bqF+LnQgTgEIwb0fEbbxpybjgV
cQPM9itnorDZ8IpXRkJqI9RRnBQh5FJo4dAHQbBATqRCquGhFvYY1LH9oMyO2Pz2guCGiP3GhH7Y
rONAtwXNcbTyDA7C1i1lgY/2tHXpnZyRHvmyF+pv3ihycF7L98mac1BNWylqCGCKJOAQRoDyJ2N0
SysLeS+kB6BMr/IE0lzkXvDgOaO4s7nrv4fTWwh6yCepBOGJbJUHWHi4ePXW4sk3gXSXhLP5CRHn
9GgGA5YdZ0PWYrzC+YfY7acQcRVO70p+L5PeWi1e/aVlcCDwx0Wd6yj7hZVMDfZDYmfq8qBqDCu3
ztAqchsG3UMDWn6bUjEfCHMbtUqxMotCvgtpB/4dqLAHsWmW0WL0vxFQ1UpLx8Qir8MlZ0u+/aRl
jV12ZU4eDDVYcdcHiIvp+DcJZwahllOVE9Ej/MJVVeldTzKEK1IaMam1j0fq0mYjGHBkGo3B9mrm
FzDU2HLeYbK6wFXt/fzRNQMqLCSrrfZMiWnwwK7NEb+T09O4gkMLzSjTT8v13/hdcjTvcnqr2wf0
7JIj5mmWrQnqtc+dm7jr9f6eUbk7METtqYMduEYsh10Em961rNsBtqa8hyz2+IIcdXDzsBADvwSp
v+Fnelf0OjomdEd3K0We0zJq5WV8echydHyzksJWNFlKn8ddABKWRv67pBfrXNUp2meAM6IEwPKF
LldcOoZiCt6IsM6VOu419qmZIqubh24q9Es93JemIomKFi9C9Jkbd7gZrEsU1MSSP7IaPDhVu8KO
Y3xo4pTduP7vZ3dNJ0K9bMZhgPilxNyHrVKOd7iFHV14riDli7vSZJDDiE532r6euj/dKHK8qx6F
bkeZVdAfT33KeBPVpSOjr3ccEvoNwFNKwlluqlCIGxAAvYugKeUs6nq9pnwFqdkR7SO9taMylG8l
pwLeuqsYAWJeGQTsvRZYc3atTQR5mNhHf1MmWtSWQQAxKmfbL9Ps2OlytHYQ538Cty9U76jZNQPu
eKFWBfItrUrUK/EjX5tMPx07aOstzEPoanFXo54ei+n21N1uJcDxMEwqbzzaxmE1OlmB1iRFP/X3
l84TnJV4dlPjYLUkKhR5wFJEWzPmg94m8ciuRYe+AcMChfzSJWp4WkA+xLx0hhoJCjW3bNTympVp
MKzRJ5RJxQMIAjS2HNjpo7WkkwucF88Jk3ksIQ3UGisKRwavvysEW8U9uiMJizzd9mBwvnw+s5Wd
D0Siy6qYpzwn2/TekZXFxN9ycra/B/CYzsyCY9SnatztLwjv6mChvAALZvq45JhXGiPmz7z+VF8u
ApfO1pcIbisQ6DK0cnIyGHns9832ABEX8F0S2ZagyjSQsz3rWTycjwofqqE6a/b4H8fm0SyuVqlL
XmOUnrSZNP8jj5x+afBEIslwYZILgcI7j0fYUmod5DcVBDGgTgQH177WDb44qasFbMmoWYipX9P9
yLjd4wa2TqFIXOYaKthYZmzxpgjl2hPjVJEnddejUAOZGU9K7zZDpsoc+ASFsl2VHQxIwf9ayd14
b5koCkBQxVAn7I2goiyYHo8J/N6XEahvVgFc7UCvvpCtBKdZo64b82B6D5cy+DCIawWxQwRaCkN7
DzF1GlSdMHvVyuniKuxm0jFTMyMGWa7E+DlBZ8wpLlgH5aSITs9JI0NPbLddRyN2pk8x+oFHe9zJ
/5cLv3j+mu1VBKbDlurEWxjd8sWWlgtO+xkGLeRR2G2syDeVDZFTSyVXcuBd6sf1Q4Yz+/wFT5qU
8orPSIndEAUwFWTVmxAS5onwWphg/wP41agF1Y5Ed7GEdKACUm4sY9zY0p545R+WdnviWJu4p0kz
4blxNhAz5VxLDOYIVgM/Eq026NzDqf73EICPj6TSZmd9s9dLQG7hckoo8hV3O9/eAgXR9omewIoo
gXwDv/xWR9n8pVzoTcpeLOplqHMl2Yzp1vmu+BYnA72FzwaaEehM2SUX5W2iOrOP0O/92SZpOUw/
o9PIHK35maqtpjYX53L0IaZPSjbKDTP+Rxs7e6YK/c/Ie4Crfo22h1f9tacQHEPCTfYNfixpYgws
5RkNULp2Qv31a/1M/ac6oikhZikQFeyq9mGmA7iRD1uOF9huVJoyCyoJ02BxGCVM+ZIeQhPDKo2p
Lm1zdEIdltVSB+poeQSN2+Mqu53wXCM8TZCM2lFoCLPAVJE8UJoP+tp8YHexI479atFScRDyfXHb
RsL64FiAhJKBGiB9qT36yUE67CCvDmhjpyeq1OBwE+mMOVYbq+zbd2yoD0CiYst/EhW4vzyVSOrk
43ogBPj87A49J6Z3XJKwmyjtPeLH80CR/3sU2J4kUYT3Ebfei+aZMqkemvwBbJwJA8p7in2oJa70
M+VGHwGuUG0vZitxNll/r7oYcUDPNgzSzIYhb7SMSgUnthErSXskQrqekZFliXaVlpDfg27/7dWG
SsjKvfX8RZ0r8mBG24EAEIYgyNVFQE66Qf38PXKP32qTUwR/SdOKVOdpIk/Vt2WRiUEJiALd2psd
Mw0wU2I+K7o7XsC/MU0JCWBxVKYR66B5PDmHliEBKM4QAnMyBsJYPuv0C8TeD3qhWA7LhJ3GxUnJ
hBptbmqrKlFSfGplhiW8yzt7LchupZwWYEcGTdZZwAIGLOTK1pn7YrXhGZJYZw2ssOdSRmY9g624
xRWnyfxJYQjBT82ZacqZvr/NWD3afSO7W0DUjKAoyMMrA1E90f7gYDEVvYLskGems7mQCg3PHmLp
Ynwjh671BJJSbEo72dU5AQwxmAZQfWetA2G2T16afzNHX8Vv3eoPbheyx1eBMqb9m+tlj8gI9DzW
h7fa6zojjy6WMj4F7nyz7f3YLM/qq7fK4Vz04Bgcfm2WZ0dGxgwUoqhkqrL+9fRWlB6C//eTrc4Y
92luRMzHxGrjic6D703MBOhmxx44w1XGSuk8ONUTKPyXjhSD+49rdlOnp40ra9A14x7zuv1+1AK0
gDIiwdda+hsGHVCMhoCOr6kPFwzS9zodDlxxJWlQMC3Pg35vGcauOkcdLCkPzzJZPRHgm75Yc3xF
fa5AdrhTwiWtuxkOcpzSfK0AmU0Lv7RrsA0cDoF5ch4liN0zZAZJmAafP0eBh/Fc697K8+dAG1cJ
1NCGKB3zMb/VMbyu6ySdFljr0uZdum/kNFQ83spIOdfD1/chCjrZp/+X20ngpY3TmiBeDVrbvfK8
AbaoxcYQBLV+IHw28S+So9VG8DMHtx5WDPWiJu3PX0uW3brLMbhmJucRGZlKOlkyoLBDfj4GceLh
e7K1IAh+ia7jgPeUh38wYSnQwhE5uqAzRQxP9saG4NVRINteoB/LT1jq+YDj5CxLvtBhcEgQYhgk
PK+uA2kt4teSxiZXpsWXt6mXuPOi9Q1uwrmULV76efNkIIK0AJg3nrpg3LMCO47/vL28nxspjaKi
htvAXQfp57g9cSvd/ExkBD6f0S0Y/xobnGS+dU77Huh+1CK/Y5dzUEnUp5Ma0gOS3xwcFkNsFsgc
4sAejoX9cPtlEIdFkNVdX/bdQbkE7X7VwDihY0Cbc+ag9A9LH8dn9oGUh0iEX5AfS+1wpleI/03i
JP4fjO7FJDFBnZ2V1VyLf+8jMk8OxK3xPlVBvso70mW4ujPTLH+bD2R2AETnFiEl1FDs3JGojsUy
IeTPabjT4/mYozf5sFBiXuB7HYFgLybiuFGKY9Wktx4rdIYC8nQvGVaCwPKBbRTV+BZZVYCPJWH8
LHtqxl1TeW8ngMtxJxEz31WmDlDbtCdEIzaQyRCx0yUq9fjUQEGK4zNbz3ERHmSY/28w+Np/Xc3v
v/Z07/9ams4vdYJM+llDVKQhV24IQPZxUSts+dPgKKxHPQGxsmObV8FhvsB6bW74I0hlqaeSKRa2
GECT7HyXtC/9xEC350y5cU3k3rkC/f/N/vNLOSp0v15UV8aIr3WxKEY70u2F9NgUa2GnFSYsUxbb
0uQleymej/lulCaQfz8/rHB17Y1Uhr0XFuSXd+5tjeqSalVMvNUdfPZUDd5G3rqOcRI11XoWeh1n
UelRswP2IwYCaFXWiT+HQlZptQFR4M1PJ6HdaFaZosmpvezCgdsXR76hKxhtiFicDaQsKg9Amapw
WmFz7rp9BSVw8+7qT0JERWA+Bw3XFFQe5XE9negVlFvcsPKaALdeUWKdILPed4UXl3WH1RaMmD85
GfXgEfu4HOan98SpcN8+kWNmIrL7orTMPOMx5sqpQo4SatNYoapmYCqAN8XVg2z4+pNhgHquF3i6
iPvr1VTJtFNO37QbrMUIXt8lhpqAnvZhn0K5pP9OD4QSo5ECpyFvr7By9/76h7qdxIzaI+1N52g8
8EQzo4aBLhAenxNjyOavtrcWL8sPW62aOCJS/BiuEGCHJdlz0tzKKPw1DinY5suDhQh8A9Xjn5ZV
yRodVvnPe4nbIO1wWyDHzhUqq+VBFa94h+78eSuRArt/xccfKTnJeGJytW4HaVj5/EgC0ilb75cz
kQFiebiKeRTmsUGcmHCkOQgL0bcbuMmL6P1dyXd8UU2U8DhOQNfA8uPe8Usz9lvNWo8KwiFwC74U
1oPU5fgjyr3odtXs2/Y0i7YJcL7aw+IfXWX+pcujox3yieJVnw/eCtkb16eQO7q7zQGoXQT1NRvz
3dGzZc130KEIoygBf3cCKioDY7Foop3iTV2xSL4tUkIUUXSpYSxluZgil54PUkjwgnWyxyp1sH7U
FvLlbSsVjlias3Ix88c4JNMd1ILtYRiSKvGxzt3KBNNwgEQc1dsI4So5K4/5vdQ/ITcZjaTRZvQT
Ik7CJFsZF9kVg7FRyR/I3ywetDy2uSSDrt1eyK7HfrmTnsOpzs7NjUGRHp7PJs5cLSTaoBWx8gQy
IgBvFoXIPRdTQ1dNokwZiZOFNpq95TdvsoJBmc80g3Rf9S8kefuzvTBUW19ucYnEmZyVKkNrPXxH
R384gA0q8Jown1cvG07lOxUaA/7w9fPnMt+5RnCHESyBg3cNqazHw84RSOldSZzZ7adRrBckE/Ho
3xW21R3gQhVn/z1xKtI+aMI7ZtJUv81U+ntnP+DJUBNAcQgbGvj76uOv2zdxQaOlE6m/oyg6ZD/o
odNb630VQJ9lv+Xx4fNHKTyHy8HgDo7UIh7A3ZfJRx0yWOlR5qae3VFXkffjiFnTQ9CwQhAdXYja
tEchtCQ7AT3ha3BgtwF0zPSunBQZAMwrfhswUbIfbv5IsE/dOzt8aHCaxOU7nSsAaYR0sG4wVrL0
1MKbjKoM+LaBwvYaQsHFFrgv0SWurqLIxJa/8JbVQ1PjZe3z1j65oRm5OaLGThGkq/DYeFrKIB/s
i5YOoMTogiWsRVPH4MAN9yaZ1yOJCzNcOTxrhSi3zvAplmN2EBMOg/ByNWJGs6gOUtza29GgtMYj
TNk68O2oZ0anJo127Z64arR4UTGRdQ+BfTatVhvzjC32QkzX8U3SVqJ7Nxq0WtoZDHJiJ08SF/73
UcZYnQiVRfOI0H8FDkJXnDg8O3GRlhVwPrV2Tum3rtI37vF15kbHOWMPNtDt69YkfEtNVg/1GI5p
h263IW298eJG6DdJUKLq/j/Hw2cA6fr2zqG+Dn6opU2LmVQcsznrFCc2vbjq8sd/Z55dggBdW8gJ
tUonx1zJ+vhBwoUw/zVkLMqMBiz5QMvZdyryO05TbHEtyMBetkicxOiqcE9NXrUWj/s8j4SBnvtv
dLroB/OQ7wz1lLR1RGR3cwUQSS9+0m1DrlIWQRauNcuAqR04qVROQpmeSGYtRAFBDe6D+KilPKpu
Sj/8Z38tR5ri0Pp+QKRL1q2rdoKuqPEbYS2Db4SST1YIqqKdMi14cojhbLnHipqaMWUrJHH/zg+N
SKhfCN8PYo3ByOpbg2e/Ty9+unkG1/5Vd+QIyXCcbOa9F8oDdxrEuzs1Yj5qTjXl2Z/l8twOM7JI
AQ4O1XyycLnYAiILPOvWoNNc0srj4JnVdLJ9QBP3xPOej9Xqv4KshBl8sCdHARgvYIbxTu5udhYr
6ZAHb0MJjuKFRgmegDrmXf3jX2CvLOGfzvrQAjLd17+qo4PwSMvo5Lbqx5UryIeSGhYPp/PLbEU9
8GpZdgEM+IGYhLWYWTg3s9HeIBH3vvVKGr4aAyauTmCZXtFhbBEoHPa439zgd0cOuHBar5ML9LUM
S1kUFxJabj2tC2Zb1tRPmu4MqiwxXc9OoMqBVYZDlOwBcsIB+QlArm+sYoD0jindale4maQFqyaL
boULsaeLdnkMYjuXvZc23ZhnOiAiZIhXxZhEiXRXRlXADN/5R7S8gmrP1GKAQw2Qcq6wTssIwPnY
upiLYrVqs6Vp9t+PpO7cSmTJdm25peKr/qGlUyvRwGyotOzrNDOtmEImpDZZUDawzYxtIlzQ9HkD
zFbUAzAyY6ATJMh+KF2RpRh8VeH7rNkqSOqGcBzipuytVHoxIX5ccGnpuM9grF7QuLXGVO/osHqU
EMoaBJ/CvXizDcnK78hr4XFLyjj+gmt+LUlnSy8Ih+ftAuyqHbmAaMptsZUCCulMq2ZRS45qNTjr
dy4IE61rQvs0Nx5GSFl2gbDsC1fwKtJKZecHXxPMkCC0zzcDSUswhyd0GZxGFtxBkTz8Bpz2K+AL
aghE+K4XM7SIOCf4huaoD3BPgJa2r18U8yjBf2iBgaSAbiRjk9jtN07pCejxas1Gexedm5SH2V7M
6hKFNE8HMjV4SuGAHTlgk1mK8dX+NpPE19ntFzf1Ss3sZzwpi+e8+YC9c4mLvNq1g49naPtu0AsJ
27OUj8riVVC3dFW9rimSjqPsUmHJSTjtxeQq0LEC6BQLLk5uxFDnYqR8v34fPd6jONSB+rf44Vfa
9AAH3zXSCr2oE3nWuP9aEMPd0/oWVHUmTrxC9TVJc4ZZJSop5oxfIAuRo8CrWwlLpRFZxLLpsFbG
+c+re7H6zIlBvmZorBNHSoDHbjZDBBwjAVLil/QBjPbwHoLTpnS6tUgpD1DNOCCwapM9m3O0/aY4
SP4te5zGFFA8IcJufb+uhvoC+tcvtGECeTe8XeknyPbXJChCESrP/N7sleaX/pOks3qCS4ciT4et
SMZQoOykjLUn7Pkxr4lVoTILNKyVyU/cuP0n3I53s16P8TF6Cguv1LPkJpUpjc6lz5VV4yc5tMvA
IuzJobK5VhZcuC8URxkZKGAU/f3NNRhveKf/DDGj8Lh9TRwpXOw/U8D7ggVtM2l3bzwWAG/wWi1z
lW6xgSEhxpfJ69ioag+EvHBcOz67+qawyN26SqoXEBE4BcXFvhRjp8cp8FH2WoBqlsQtR+eka8xO
AlTiP1EhXXyCI6CVvpNF67tW+f657/VG1SOcwBW1KhZN3985NeYHhKgKe56IXOwmMsdOTgHIrjxC
lNviJBTwybmyDbaQoTr8xZlUbtLUaYpRgD8xwDDaaExmaOPH3zLNnKOr8b29kntpoj1dNiKguVfv
5HL9Iid1UB5gl7Vd4C5ekyRXF/HoPJnbG17XhbZ8TJD7wZNul9VcTl+cpt6n/mIo+cMtEHjEhZuM
1w7d6AFh6ujmCb92en4h2Jx8AoTlkpGU83kZKKBkx7wQDZhnAuKsNRVIwPEO2bJVgkSJLnijrkFj
msUptfxWbjOa16YFQiCZ0iAc5MY14XAFtgg33VNyKakNIdM2LIsanUTywkXfwRmKRM1LNjyl65KW
BKIDb6Iw3YL6VqdyILI2kPSH3TsqY9N/YQsiCGdTJrV6aA4G7hOWLz7oIhdleiFBfibNToAja495
tolvUSNI4sXIk1YABwujKV3aWsaPYQuMO/9iX3PZoZunMQDT8C9U1bj4kzpocBDH97mc2rm949cH
6/ReYVUQl1e2kjTPbfLj4YpuBT9PJn+se/X/JVzR7vIvrzwhXja5dYukLIOO/qDm4gg8uSZmWmOF
+cgcozPsCGdSi6w3b5CdWUqLH4a3ZWXtA83j4I9YrHIPkjWFN6Z7wxGE74EFRK4tjMiHltVaryYe
lqzkxxIXLxJYZ1aGKnaisIwvqbTqf8qwbV3a8XKLtTzSBfm2XsNpqc2ISJnlOi7lcYsQUtCLQQmv
zo1AFkRk/FaaNBmF4RK56ipmXI4J4zbxSuapTMS38joFe8TG9seLVvGUWhULRxkE5PtoKBEnuFlV
GGlqnLspjVvH14sq6aXUuMmi/dFDxr0IEoCZe/CPquQ9xn4KQo09WOqkjuQrCnIywiB8KdeuqBOm
ZBMYbLZ4qx1UBgupJNl84tv+WfpI878J73xW75q49qyI2Xy25axrJvUT2zUfDYmsKM3H7FoASdBL
lmYbMNcLmy69VlFG988XiJb2kI6tUcB4SalJUq/gz3VjS6Ghy+/5aQGF532lVhWuebgHbKW24m3F
0rCTAQRWhePKQRX+gUPxYq0exfX/QpHYhPA6vj1JPhIjTt/K40eEVDPso0H97NMWQ6dZwhhQLSCu
T8k1RNgPhsx2yorPYuwlfmuDPEhExn3ZJE03xvNBds8HEsjsc+fIjAZkk8aldcQ1ZR+g/IZBlbNq
dU8RIhUZPxn+PDgtYbrpcTMo9i7vZmWADlP5c2EMbCzQMXsxTQZlF7OdAHIPInpNng1WVx2dRuKp
QVZ5bKE4F66GuQhNQslENDkCvwNbE84hxSMS+YrVbh47xrmZQ4mJx7Nw7awip3j2yPowulLwqrjP
7WzKRrQ+x4KQxf/HzE4m6gXCcPwNMP23cVtfJ8N/XW2JD1ZHyPCwojh4wJWnlQbZpe+PGPSHrH2a
vRWkMPNFxogLVIVcclxjSe0tMFZt2j+jdjikhakCWIrWYcy1vsD5l3cE2BjGVfMFVqmqvM57iUzR
eJNGl1QYP88dQUsLk3MJd45YGVSPtNneZ6y78rtgzhBWZOjCw9b34Vhi1QlxRcJlHDEDeNtkouSj
lr7XkwUq/zSNrShvgZxP1Dgw8N6qrMwYh8Cvq3ehcPGk/LymNxbNnHLifJM6S7Xlx+kY74Lj/vBg
JTA98KXOiR9tCu1+BnkTduxQkaCmGy4NyrPrT3kOD6VuaeTV6vLjuhbACOGU6HMPtbmdopjA8qjv
plzkIPkfpv2TzppP5ImQtmu15w5EcHMK3J32bklQH7Bu8aQcKQ4IiiIGd+vTMDsTzjflMaiB6RiD
Y7WnFBQccKa/JmWN0Eojj03wL7f23Vbn0wB56/PEkcYXSzhbhDBeoQje8NyCz+jE1g9pCZ26NIcx
lTKRd0scyM3auKTxTXF+taU/I8DNhUr7J5n7JE5Dopvg2eSZud/0RFca7PqmhZXTDApT9abafKsV
yjt46ToeWkCmGV7B/syxbEhTRpNNbWCJ6ZEHaz3xRS1AxfLtqrR14dC1qd1+BsaGb1/yCV+jr2rc
t0ftRSBo0L0Qpj6a+fCEI5fIDzuJ36HDZKuQPTLUHlbYSdfA8D+UBWCohg9n3eyEGptgRi1dyxiz
LCJVjbLyGf2AWMlBLcT5EMoljQKqrfXMvVXcnb8bOqmj/C3DiZgELInCfhv2DDy+th+J6B3lwhWY
k8zZKtgxYTnIcqrlbe0HsqdBMCO8AZvxFG81k14hERdQPMMo20zLEERACuNhumMpVtKounHoOP72
u4iJhEMnxXXs1qtLuVHGpoFFLZsxv03pKE0DKofGx8wQqCZDr+nlHW3IKqFFjnyQ4ByVGL9x301g
l86tmwouRRdXAHlrGAlvis5VXCWkIQjBPG/FSVVapEKEIjhHWz/Xf4qrW6UYvw0EFDz7oGYNnDvh
rBnZURe14jaDJVAdbp2YMBnUzIJuGfcvfcR+sVy7r+KPoa2jiYZ7ZrLXPGCWcb3NW7xpYYVcAAEl
9B2h8bI9eB69QEneeyqP5QNfASOLwLrxyemL4ah4emWBqsu72xZtUXen70w5bvxrTDO+/GrS0uH4
xpejoiBXkj9lKvUx0xYB9QvZQLJFJt/FDtw4Sc5NuMUbjRn3oV/hr538axiD9wlJPoeic4505ZJg
dMj2vbIJ15AmCalLxzQeI14TqLodLKd9kBZPKiXjbGfuE+uwV5x3464kBc+XmEWusWZXZob9bF94
RKz7ikQWuEEGoe/2CizWa/zyM/AYOpgTgJCq1WNmyGe4W+k1H+gC3/rIyn9Mf+DPB0UAkqt/NkEK
A56hUu914fknz0lJNWxFPwOtI4oicjetQp87GmnrfbbI5v5sggth392TmEmeEX4jwcWPWSoJxA8N
WRWRQ5JXOLQVHwkeJ2vfajRTwt6NVJJwPCU1Y5IfjWLf8uv9kQUoN1/yGCl3BDzSj/sZ5CBwCtEH
38gBN5PSwe1sGnSiyor42lQgpnlolRwIZvdnkzct5q0AuGyuvcHwSq1J5Vh69JvH5cn2hp5ESWdP
RZfUzQIgK/KB95D70uPpcRdGzG0vW77Bd+9jkciHsOn1UcPk5ptKWJQv0D+Q7VpXtI57W1wdN4nX
6IBFwP4a5GTi4nhcMWvQBKjahwgqSzJBnHs1Rb7KcwADiKzSDZIxh3dLVFIXnlxW9IY/Cf6FXLP7
yACzA3hVSt5h3fEaHIH1OoGHxO1oerzBUA4PEtoyitHtYzp4IG67OY5/w9RelrwCWyo1zKIi8ZAf
1GcfH6B5rshdVroNPKzxXqxMpuK9vehmB1Jh1xLv+PgUHt2tACMjugH+mXSiRIAm4aSvyX0I4m3X
CCfEjb+HzT4K2uZWwaleoHI85dqq60J+LfYMHrf9BO2wxJmS/50SKIGF0P8hm4pOmWvONGq+FUAF
YrCK4k9skDxlWGQnI6rpcDf/OR1gnsd8DNMHvo18iAhD+h2gK0VJJYLnDCXbZf5xPpiLOl8funZq
z3dUzN+g+0an73PMcz8OkS1qSle9pGLHZUcEizQFKTE3rNyZTPUL/T4R6COF5MNqeOqrWMhZkH5R
X9RBdVteWFw6nFMohjsH44N7iICswaunpa7MPv1h5byTw6RFTb2yu45Mh2myGm0qR2CUwvJ4io7E
CqU5xcuVLrXpCkcUg4oxOoGqvGPlI1LbmERCPenNhsXnGUavztpyUJzRgvu5b00gimhFr0vKJBeM
YjaPEdxDGH9SHJZ0qZlMuOFoxMBPucRv87IUMKrtX8vMHXSOfjcYDHwOQ6tDOyikpiIC0AlH0ogu
g/JXmKAcSEKc4hP+8bhAVwMVMsc99BFevJR7DI8rXBSrODnB4RsY8ydZJmP8JzgXqPNm3H/sZFhN
2nSzyJH4Vzv84+v0oxbXXltbNAepJ3Gi3ibkvojIEaJiWY34OJHko9dsMX45DLhxbIItgeIW6BE1
ubkTGEYYrg6pCoSWoE3BwA8/ZLvnaXc/eL2gddkg7nIAcl8+veJacvdIAjZUX2F5J0G8n0N63eFL
zZFfrrveN67/MP4PTcz9gGrxTIiwRMX35hC6RjVOOedKxkHlLIFupAuqHW2Nl/FEdUH8TOXuUo1j
jCyLVxeIDX749GdyygdZFH/0EQZ/2PzdaLdTQHuDaFzhM/E+2xMSGmM2tEFACcKKE4A2Wx/Vna8l
vDZkgHip2YH+rOfSuOMC5jschnHWneyL3XZEy8fl6eqcYOKAXv6jPxWyGQgW6TMQY7dub8hm0qop
JD4jOk2sZMpA5tFyWAsfvmINSKz+S/tAYuxnauO7KqmWpX/kGsZkSZkxIs7tBgKbhBRENHg9wxQK
KZJV8Xhk+7g3pE51m3NQ2wuv5ccdkE0hjiW6uftGBVuLcBR0o2JxGTiLoxKAuzYTTHXKUGHNhd0H
v3+sgl/wkzxRPRRHWxoXKM2iTjbHNCMZ/LPXsXk0Dag12W7ZhWISgeZMNNO3IxMpXetZ9E3XdWrZ
6JL/Rhc6N/cCd5pDeAls6NM5Tkjwm1b2KvhBLHwwCWJawL3DHOVBFR0NP7ypri7x1uavAvUELyMB
yeWS7cglP1YK7msP9Svx9CqjpRcJyHSWzOdXQdF7jk2e9GgJrDQGF1IWHbnu+Q4kYnXszshGp7Tk
vcuylOuLYb1FNYUQ6MIAllJxix0mtNWfpHC4AIehaEd3EmA198mSapCbPcm9ATcD14kSnYgBxYbn
Ibx8otfZYhgLZCxKs20WkV3Hkgz1To4KkxN2KTOKnbJZCvYWwGcsRSISlz0HbKXPSvMW6VMtialS
rGswKNHv1mV/Q5+mcqNZ45YI8DSmFgK7QF+Shcw/LL/7DirJxPOpBQ/vO7Nkh1tSRghoBUhWB+K1
REYe8hoSuEpsozcqKDEDx0yoCNnTWH9Mlf+gzvR31td6ZZoTiWOuGiCHgO8975cemZ/mDNtsBhDi
SFJ46ngCgwvToKgOdmEWEQ2oUlLnC6QIwSIdLYyjxLDZ99Qugmk6BbqW1dvEGwjZdxOMAecaphk9
CNMffSeaAjKm+DhKeM0N/4W8KEi6bri4R5DjUx0ZtauMoviOYggeE4KZ5xLXqWUERz6tgLLuDHf2
MobHV85bdmKeTruVl0TrJ/cJbxL2nW6VaimLsA0Ext6UOIArC7BP7vVCBkzOl/FcHMREdT7KW7yg
SqmNP54ncuuUN8G9BCooLhZcL3c9s5DdXn1XBcTcoRdzYZEAU3szoTV1IZ/u5dogP1Mm5UQ3+MZx
zq3L59NRNoCOqg4uLeRWXANJfPcIiF90fw23oaqeo/eOYKnKUVD4BxdAbPWACTDnxqgPMgbyI3bx
s6+orbrvQjo86L7VLQut0DBsopiEL+yoUp+FP/IflL8SVNjxh9Ug51gFLNdP1FkTK1ORbNCUEu4y
LKnLb+sUp3pcNDG4KHvaXi3ryx0UfhAu0PI7a8BbHqWfz9iGsuaK5zvDgE6YwjwhWGq+Wwga18l6
ORrRcDHMqBVO66bOW6kVLFSXhnt0oDUuw9XAvn7nruWj2U20s438FXvuUCVrRtCJ8buAeqlL6g7h
iUwbm53/7+YjbHTuRnBXBJgiA3SW7N4EMhPIfPXqm1tl17WyqTqPPF8C0ivfJnmadPqjGd/EJXD5
ly5jLSUuequ9Xz8XI+SW+eKc5jxY5qg1zclg3w4bImvY7Oy1FB+ii2kxMbyGFYeZ4hnyYsFNGxVX
/HAggAmBvcR+y0nVKKCLU/dwr/6tbeL8XFZAmtwGlkZo5tRkNrfXaLbtpq2RvNNaO8uVypOQ7C+N
RjgNh8XptI9+SuixWigaAejj8dVRwOQE1K12fkn3eVX7TtpckhWB5qNxv0gIVaH5KhLjNsFreJQc
6z8GLEufMeoesXFCCCe39PbylbqHv3mYGmVbm63CFkt3cqfs7AUFa/xZqks5MK/vBiNl5GCIVckf
2kpbj/oTGz3Rh1pdJ7FRZg6mQ1WAz9P89Mj2Pr8ltPBQ4JHy5drPMaEJ0Pd6JS/hL1oCzdCvXhAF
/IU5u+CXUx9m3pEBod5JS3FJCIYHUGJvhb2ERM5Dx2vAfrnhBP/BcIxPV6NuREakMEWOyaYDw+KI
FXg82uZ8Wqp4sb+jcCeCMHW2s9JS2bvCYhPrS73bIoxMTPgUsWwoJCbo9ZpbluAkEgmTkCpOI/Hx
NTWUSuXMq93iumE0FsXDsIPcreATnAmvdqaxa8I9gM7gwWUXobNa2lFjaodw8RtmvT3O+ELZNvT6
kHSSKYd0K358rspr5V02OAO4FZbREgBa+dle63fwxGCPAqcn6AeUG/G4OaGSjVQ1ooBfbFmC8Tk2
BxDW2xALnuOzBEay6jZ2SBGSLtK6itDhXh8Z6puVGQ6LMsx8g7avD9viHRNUnbsJDe2vax/hlOIK
GMdgmAMvUTCyUt8tcdOhwwAKV04dnHf+DfocXu6+g0Q0Bon5S9GX4jw5FC4q6oueRZym3aX+RHk9
dTgsIjfPpr14jgq888fILbE4I2p4swEREiEf3F1vhzYPhDM1khTseXZgF1Kdyu8TNYs9bHIlIgYm
s5Ui6Nhv8hCRqgJqRZH4qroyF6JArYs/k7RLzqPY0/TYYszKG0wdOuwY1kptJNvnfsFRI581c2so
Mirkr3KSkrFEQpYA6puWhSOOTIYMcujH1WY53w1GyYK1AS1yw0i+9fkr2cirEUHaMElElt/FdGzM
b6J+WoLxKDC+UkcM/DthYcdk+9/zoz40XRdR1NEb2GzjYXRgX7Gjuz/wqQ3M+o/hns+W2WhYtyoj
O52drJAaEPNfUnB/sBXu6voQxH61bTul7HoQT6yPaROtJIcF+ywqW5gd+3kM/nMglbCudnldtelN
Z5b/pCMppmacRT7rsK8zl2PoeUNFVjLGW2uay04AFA4vbtNsQUv83vnylbZrADBgH5S1B+Iv79Xn
NBbgVgkd5WANJO5sV96iykl5ecVX9DfQAG+AA6wZzCShnUNOx0TeT89Cyl2LC9raomPk+Y7hho4A
ibHp+FLZc0X6WpzSEJAwGrNnBOJ1RJiv22EfeAgT5CpR5UUsklAkiw6auCZbyZt8GClJvL1OQl76
qz3vw9Ih/LZow4udU4CDExlAibVyec/QiKKEciGPldaP9iRA7GEKP/oQpnLs/M42KxW5f/EVdnua
D7wb7uRiWuy69qKjG/YNTdRpt2OCzg3v4dnHhRba2U6UkaVK1Sl+xtYNwli4xiNMTUfDgOCm5FNQ
M4s42wyrsoK3yh3KZd+VQ7bZ0ay7fgqLSu81zQNI9AK2S0vYWr86VsOuxXZcpQrBd6OzVM8An9dV
8jRjb26Ss+uT4i7+DuQG9zg8jnCR7j1EkeycYwmskzLHmldP3xRMmdEFu1b0faiT/rYVlCBNlp+H
ILIZgmJgwXJ5QVMAg8Bd+JVBpmCMX25V1jhvfWTkiGSpcl8Roh87AWfXcJTjPikkmLlxac+JXvLX
Uqk59ISEPv9/FqlUMYAkNlwruCNzrUCvlIfGivBacXhQSIHUciud6gRhXt13gIGNg9uafhHDjUEb
4Xr33drR2AOGtmHUT3FU8OHdmR3kYj5Rln/Cd4rEXAKdYWl9aea+LOhehuMhohG+AOgoh5IQhCbG
jy28QU5qO7vsw2mdmeOAHvpdoagOiPej6RasvotV2CUOd7GyWboahXp8Xb3/fgyB5fZKv6mA10z3
/vadRnkTyTx3fpugLUh03gbmGTyWvN5eIMJDZS6iYJ+STjBb7WgY1NBLqG4xwJtGlguq6wpHwrT4
G37rAqJkdFMgVhVko68BDBVSb/QoiVmM2sHK2o6e50dIeD3vy/S7kMyS4ZbxwOeG0Ckmc7f8cKjL
OzQKafXFtwQyIKMUO/Nm8Ze62MZWCFajzp4rfl0M1KHmhHI7pssx4Vcu2Jf/eZ8SyaWxuw0Pr3Ka
C7100vB3MIs0TnjTfo/6AmVgFXfqs3SU9GjSVqbuSyphR7I++miuUUNvfxxyxpXK8TxLxvspfDc8
k4RwHkX0SMZLLnU28/jC8RL9UAV4QRypiCYLTyWv4C7YifXHptCr+eIlLG6U2oSmQUUkKRN1hTBk
DsgAdqGSWBfB07GnTQZHuSOaR+t89z20tVfl2oeHVYVj77OZcYsqMkYYmdeWasmJKh9yW6Ub8QpB
qjgrc/MWbjqeTB4XBTMKT5McEYg+hPVjPZN1oEcXcSXJHjSSY36JQ+mD6ijo3D6lueNrKmaRKOzS
Yt2A6bFRI6I0TX3+0lWpo6AtQZPQP8AevJxgZkeCX0Pa5rn+/fAa+WpFgdwY4ttvSVh1qYaQRnB2
mUBUP/eKiO4bgJ7Fs64H5Ft99xWaQG5BI9bczbBbGTeDm1f4uqf//WpGHLG8iiMjreVAG0L0x/hz
4Fy6Rpz786pQmfOHPNGmFaLFAXFMeHMOAdJtILeT0tCvrpBS/r9W6iVKi8qydZDVSbwya6MZYGBv
/3FH4nOP1EenDAiUJcEI04kHArH+3HDq2uaTMuEXgq53BF4HiUdP+yRNJ4JLuDmB7JAvwy6NSgE2
aNfNzdoEwRYr7qkga3L5KqgEry108+6w1rCCmhRNxQaz67IOprWkJDlPqpUkVJwPmlGbkjkNgqV/
lHcYFth1ZRJ7Cw4EryTq2EqHROJFtqzlSTZNQWRca6MfeiEzvEAHM0X1eZaK0H1+rpVh/RCqwi6S
MKdbGa8j1k0VLB6rGR4WefuzlfARZTaAsKiusnVCGB9a6DEdAHC7YagZC7zCarQh7/fU2SoHkv/F
zKnLhbt6r10MHi/MfgHg36oMoRODTgjj1fmW7PgBnJ/hHqcjeMKhyxDYdZ9gkjeUTgJ27GFmgRKm
VnEH38Q/Qm72dU7ljlsW5Ktrx2pCjT8KVxZd1SnCIHKx6Pm3VV3UkVjt6Ua5I6hJ1KJ8zLKr4JRs
u9vxxQk6apivx+3/Z9PYmT0w9QhDwDCBDkXYqydPU5KoRhw2SMUOavQpUmewqFdgnGTQAzZuKqqm
k1UGhWdWCepiIzALaIeWz6T7McwiLgpVuyPRiDt40Jzkmf3HD1xq7jTfRh8v55ZS3J0aaNsMIisd
fskCEinhAS4+e5t0wgTjtfYqPWzplkauGFp8n/VPkinrQucMcJp29OaQ4TSaufgDRJZs0ZkBPG1S
4uShGQG+QWl3MNbhfuT/2MqF5XT7A+8srp/7v/dY8HCCC0v58l8wFM86E37n0gsl7SVhGrdq6xkR
BGKC9Cm4VVZLF2I46iis5PD03EeHWLWvxoizG7f1rCXQ6zOPOwA8JOSXejqtmylNWtVcUShUnLWl
99aJP1KKt6/nfTnx4Sc4a6P+pY3jyThUo37G4hfytu/QKvgGAmVB8AGl4dBPnwU6zOVACYb5ixna
yxesAaQUSXxAvOhpgcMw+oJDt3unYBbvg+iPC6jffqpRWXObXcd2f912h1/FE2Q1d3fdCKMK40bz
SoBVkXvng5PA5hQNO8b/5akKVpYp1KYB1//TJWPG3CqcbhVybtL1VI+yPGa9XPjdbSQBsx9klZjC
VVhWgzn7urSLBUbcrNqB2fUTC4n0f/NoMvh3VRyfLIQOkvoML2PozQ12NdpBy0Z1s4qR2rVhp5Fv
1aCa8361YVVAktST53VY0FvA7nW4Jzm/XrvoNf+HUHBynDMY5I5jdA6sZFKsGioxgfOrEqZoWPVL
Gm2ap5ZyL8JAQnUUz8tlmazNYz5ynUfXD0LUvL6vcWyloSfFreAShos7XMfvf0P4AxDe1djNXyK1
mO+60keUXnkCznuqz027gyeKe3yfFHQgdzi7bcW+zsQ35zv8LR1zkMkV7GYPTvt1l/U4hVUph0ww
ZWOToXOKCedoYXlcoKbiMisBp22/ypsMSa88ZoaA/gtqs0LvAO1AwOqXLbLtL7+EDGeTwOY37ECV
obH78DqTPGUqQ4cZvODwjHvLXQWPDgyAf04W7Z8XTEobcaH6YaW7VgGMvKkTr2Tv4HF283A59roX
RcLyWwxhwchGfQEDNvLkijZXFgV3ZdbeTzimoDeh0gJSDcRdTjRrOELbz09NRHKDZncGpPaBJqBd
E/7NCCL+1eTbZvahNOSsrRJerFkJ9lv9878prcWrCxwlsb8CyC5717UtcA9eHhC/MxfnN0dU8dxs
llHZEHmPsFI1nx5jpxq4pRPgl+3iXRVCLfEODOe6/6XnWT0f4pOixTinF4wsvm/193tr4vNGCjwz
VqQ9NCBMUTgcbAG91Y2YoIGTBz1xzvsryVyqAFVqh8dt+ACHgQnTTTlLTp63t7FMdndScKxnQfnh
Z2BKBSd4SA44kKEMNAzDAILhpwFLitQEibKwD9HNDLNZcWKQvOBJM3LLzfxuo7QOxqzV1JEi+6Rn
ycW56VzcLuRBreQLGLDTXMz45Ocvj5i8Vj19ss7Pp34zH44OiQZ4CF6pJ2Ba5hGv0xveLIsfySG8
JO7rzVftR4SoPuKdtHSRwKgs5U4C1978NdRrwMf5GUxLrxC/uk68QG3dohYyDw/5WO3cpe0kYaOz
VIym9GHypa38eXyof1FV2mmJeC9mdZN3zW//q8KNIBcI2bl+9z6bq/JdubETHWanghSdmf01YRxb
cVEhsefSnrRokZYEBJ4EnRmE2MXnZDBQFSkB/SaSQ8spM8eAjJjKMXxTQU2l0RSi9/dHjlYd+ztx
rRPgqOHTfqWZKP78CdSJr7MNHvt6UoMW8vMKyzHMTDEi5DllN8YK0SJR0YWCcISGaZyDF2Jk91pr
XHVAfVEobDjsd2XzdZrKubRu3bTkps1eemjzU46Tujxi61eod6fZG8h9bgo8fJHb3JgTonFtXTOI
sWir5L9GditU1GS0MeBVvfwbsafbuaE0vfdqXhX/RD4n+Sbc5a3a0w4pcB0ume8sKrF77fplu+OK
g4TNLrcr4cyg6XY4eAWw1ZehWnZ1x/qdlGdWg2AiM6a+QVaL5MgXWSuNfXfJH6PcLSvFl0tE2rP9
fJPiRuhZpkZwDAQmKbzIEHNTCuden05AifAt87yZZDmNx33eR2c8P07AYZLkgzz1CQp2+H542HD/
J7R93vBa/eDcNrmkHKRpQzouuy0hEvc1aHzQcP9aLHyszn4PpyRcBIgpeXojT5knb+sA7hszK5sP
e9gmqjWDll5Ipixwn48eIfDJCCIaXh6NsLVHEMW5rPK7K0wns8b/aGVKk1H778mTZpxS2iQ312tV
0S7rOPiplg6Ybn/hCmiH4VdC10wHcHk94VM/uNctvdSjx66+mFuK1a+eWi68LZuKi/axyH4ZMWGO
oqmcuTW9LNwzHB2xHQY40Drygtoky7zu34yKN+IY5xdK995CHQx+PDaxMoVO3tucUiJRQtqElQgC
zsIALR1GBOSm0SWO7EQghbnlfvLJDSbdgY8TcMtM+Bp50ku0lziyf8nQauGiON4Ch6+PitRTzTwk
ADoTo8iZa68KS9ut8fqEnQhKhyAfcIsDnugZu6BE5Pu3esegsX6h2yeIrreerqFGrQtiRGPPbT48
pF63b46Sd32rbYXW/5gTs43UsUdfjDij+doNyS4EL5aha3bb5omDh9lXkbbunUfoPUy5urxAnttH
/jffUO9wvFgxzFkXK4C/4VbbMwuX/1W/o5vKx/ZCC8jZkuJhiZEz0APmLztB7Yq+1y5px2ey7ca9
HQKp/9///uPMcZmh550HXJgW1ie8nElaUBaA8x/0zOjyC1EWPwRZePe3v2CqZbPL496qIGv0530+
oKG6lDQVfJ534c8cV9LK4fN5a02wPW1WF40qQSWcAhHUv7BAi7qT18QobkkO9o5itD4Xpt45NLYh
4v+W48ZCHa1UTJWR0mygITEX8CqZnsLH+WrVDj/1Y4x4aqLC5sLjYp2KSIrc0PWuLyE31ZOP5qsm
GC5M8eJE1JeBgDZXiTe+ZnvDDeQLcJqOW30EImrwa2i1ZRAhY2mq4CuKjgSRQLDJ46BY25pvNQMY
d8GnYRRXhUpi3AeBET59ozNvKx2LPVjr6u6m8SOr91W5sb0ieHQGUuO2GVY/NI4EltGf3tz9pEP4
F/cB05i1NizNa6KYEWop8X08oY499V0+lbgbkeGbndr4OiabRiUGIWcKX8suvolnu3cS4OZHnuzB
WOgk1z9SE80eyS9aoaPLUbNoXILMHfC46CptGQwgNN4sI6ikOFDgENyuZCeDuUR8UuDuCBCgt0Na
ZH/r1yLzm7O5WUGh501f3IhAXJ4eqKSltstMGOdcqotVV6AzKCZx5MqRDmL71bw5hOSaNSQCBFgz
VaDhO1u9Tp2c0Z3Pf8o/8e4ldqscf7dAaWGG8ZRPtjZ5oPT9lA2vy56T5kNp4Yf+2c7s/JYrAchd
pKkdhDuBRMY47q1FPncPsaIhg65efeoJVQy/zXwHI3+iRQkGd8Y8eX6h0sO6HRMVJ1/rS1Nh4UQ4
4MpO9mKjpSD5IXZuChrkGNb+lD9J7y4I6/0E1R8mrP++7I2TuLANZb/MiP8ppFl1699N3jT+bUJb
4uNk8LMyjM+S2vMcyzXR4SmlBzEgnZUUK9wgokOsjYme9pKJpolsLCXHbCs0DhiTNL/wJaZYZmZP
rzoX7PiCceNBZCdgs7HUftms3C3V+L/0OzOR3UntXeTHP8PNg4uFnVw0ZX5xCOevg011W8U5UA7r
rvyLEaMXXxupE1pUWtr/sum9Gb4Ebxz5cFGT2slJeBckIhNQZl8vHU6IJEw+9dshwkEvn4eABJ89
MlfiiJJ9U0e1LgB0HwUKvUv5X6lRsrDMH7UBZlRgqRjb19rOYZZH67Ifql2nsscV1aK+C7ne8QDh
WiB8wkGz/hLB1MSbMp0N3ReZEjRYyeX9CThdz6NUg5wUNvybIlecAxpEOR810zwz2vvSqIrGhgqk
gitUp8t5VNiWhecEWX71GYlUDMAPUFGj0qUQjoTQi7eqTgKUUcyxSu9V3L09vLQcR7Pr/uwRa1pk
/tB8+oumYI4nZeSaxXO05SRi633D/podkTjVx5jeMklGP2jPP9ym8ky33KW7RLx7dZ7qT+LKe1p1
RJkAvvgpxq6ooWcfsutj4TKGFstCz4v3rqeOM/XTTwhGeUoE0V6zoDVDFYdzrfRKAmWPghVsaRam
n6G4UBHCM9bgMackQ/m7yvDB4biKfVIL3kH4y4dQHqoThv4wmdD/bR9s1oxRGFShqAxqghD18e7N
qyBHN/W51esygrPCKLtBEdUfCRb4Tnbj9t4B6ciRXSCLGulW8FN9lMi8LQjkzSSdGcztRJHlEnjz
jwNtCUPYqljKgMQMFrjXLAM/b4L6w65bUY3wbzac+14DJ2NBGtadZ2I4tGuPBT2P/bwmV0JAOb5Y
C75MKGn9E0VeLnoZ83qiKWksoGEjckabYVxd8BNsCxY9//IzGfR2uFtLLocQKSMLP2mvqr1ti6SY
CUwZTK3gfqH+XD6GZ+twX44MkZ901my4q6GbxTwsDljmUpkzAu/rz69uOeYE/tl7sts3F20k/mmT
4ogiW195jab7Xuri6pG3DqoqbWlWbFsK3v+z099vH19yNxuBFBN1ajFwcZCBSB6KJa635/NasnoX
S1XX6Vfo8a1VFqcLct6eoJSNVR3TicFPnGq4agYGEcdN2b1kvAaxo/mJdv36C0KtjX4a/KM5Tjfn
vgLhCunRgFNJe60Edsh7YKNvl/vBWBPUhufTN5BHQ4P63QCiifkEw7ErGg0S38a/9FKYWjtVEyob
g+TeUDcVplAIzUGWholEAhxg9fAJ3YwxPJwhW4QiAhrUFOzrekMTBTW4dDV6Vis+TT8v3yFIVwyM
OB//TCWMO9nc/qwBNIuRpZ7MUImjiduAyzbLrU4C/EypTpr1IsSdGPg2hAb5rlKMQ6qwQgd+lRU2
VBKZuXeHkUv6UsAc1wMDjloYn+3VYFP4JyZw/03oQIP/mCmVmBgoDQhLQ7Hx3YcTQ8GJ3eYInNvL
smr5fu1Wm23AugBMYhRI82XPt6YCG00I8QOVukfkpExTrNek7TOSdmF+mqP//4QW5uiThPSi4AvH
4/O8ZCwoxrHgtjkD+V6An8XtFzZzn5ovj4IcR56FDB1DDdyX2YBtciZNeJtIEF0M/AnK/VnrbVIt
pPKhpDnot7ScaBDq9q1Kcfn27ekw/PuwwBUJ1DNyXuP7Le16epcnBdCh+Uk3ZHQ+YJFovhy5+vUt
l3KO+/w9tLnAGTZFBua820PDEiw1xiqZtsgOClKoMXfN938tN8D17KeKwtHfGy0Hmvi7DhrIZJoE
cAeyr9C0Xjq5HvXH+uz90JQM8Jbu51fwGxeX3yDIY9PGmxOAiuZ2evhBWrp2j77GqUitfXH5745J
ZQvdChxztlRlElmIZbZlZW2BykX/tiabyQoTmxpb6EHG05kQI87kyTKNtaA/DfKxlOrvQy3m+skO
Pw4U2vMPXerxjMTkt5SBDS9DVq7Sx4GzTv2jEOBMhjACVLuMIO8oxPGCoVMso3BIf89VvyQrvbnt
D0/b0SMVcc3EssreybE/AYTZWgg+W5SxIavDhl7qhqf7M7tNfZaiJjK7dUKmRUIWYqd0wBvFRXx3
Gwxhie+bFLU53z85eyGdpry+rciDwz3iSyoQrYJhetJS0TwSmVvmXpDO2nkZCFupsy0bE+eMnCTO
j1fygOvP1OIfyDuCmjTd1XuZTh8lGEXdIJKb8Hz54BWDvRGHE3MtW+cD+V+/d3TWVtyZyXb40+r+
8RNw+V7NT1W8iB9Qzg0wzdwlLkMh09BLSohJxg07Jm9teYzv0vbqtS5p3olOKgcm1DGnlqhEF8t3
U/SH9xkSsPb72bHhVuI4dL4pATdtXQqStgG5H4k0UzARU/z2L+DHPBnLfmZiR5GPyUthgzu1nRUD
vz9Vr07tLgISMHD6s1I8CYnIwA9hABeY6ZbPrFDBQd3La+TMmBf0rFFnuZFnSjxx3NNo2nsI7uhR
DVNOm2QDZdCyh2WKJSM2cghwbxthgHI+d36h4mEnX4fsabOK3Bb1VOKqFUi/VwYUZVb744maDky7
dPmSrskavgtWF8Q3KLWLJHf0gxNDD38g1V979fBpnwa979pLa4RD0Z8imaYiZokTjxUuZTw9s39H
mbZdMea17TeZpepL9jl3BhVsiCJB35eBEJVLl1GnHTWc/KpJHHoTEuouMwXLpFCmju8+xo6sqGu3
WNFsXbcY2DluuslV2Ke2cHsfFWP4ZuxMuktZzwClTaz1sGAUTUH4WHGe5TKWMpZWIrBvfnKPaUEk
YW3Y/J1yWNC1zGvjeh8D9Lz49FxzmCd88NQans7Ayj6+Hyh0VTCPH9KmKMtIqd+H55K0IifjwRGA
ywJAbUIg+fkdRRYzwqeM+uawEwNuYuMo9TKv7Mvu3Gw8oUkZPVNfq5ybvBaLc31F9nO4Qi/JfyU7
U9bD9vOrlqscJvYesNpcOoedfIsf/ZmB3L+0juWJ8ywrkl57fli4ub+kRTieKFFo9gte9oQAY7W7
OkfK1lJh+D0uOilEDwjnpXwKberHtVJZF2gPuKkyqZ6z+ytdQvFFTgcyjDL4/+/5nt7/gAfRZBYN
CmfxPoqfnPa7GVVO/ihecOMALAC2bb7eStwvmtFRTSmfb13h9DZ92OrwjeGoyf42fvmeb8T6j18Y
PjP9a2GD6VAZCqMakSXvoeM3GtfkflPikjLyKGznfpbQWWKu1Gx1C0Jihd+voe8ajVc5tw2WO3UT
6aiggmN1Wo2f6x4qGu3Lj6V0MWgREuHmBD9u5RAJoq7Cqgvll5Q3BLsRUFNLlLT/j9tzAyJBYSIf
WeWu4hQwMKYbvA7lSJxKMKy0AFXq5rYaECniaNQ2osTPdaHAulbj3aXjyG4S/0bupK0PGdjC/9XC
kJ7Il/kIP1TNDGcOSWFp8XWPPWkiVxwBPnV8RA+3Vg6sxfAfivvTL6m2rEt1rGoP3OjDw35ELGq2
A8KoLKyKKFZ7P0sJob1zA7RxSkMnoevS1rW1HCSzIOXN7V1KxzaLkEls2/UCB/c9yuUXTWfD6dmT
J9B6b3YwUW7tx2f1erx7X94tXlkda6yVmrxfq4ncSJ0UVXXTLY7H/jl+xIFQWdnnnkuStl15zRbv
h0JI835+aLQuuLaCfpkXhiS/WFEr3T34rvAO9vfvivDgvgg0BnjCixZjCDXUbNlelrgT4/+10XtM
bRKSjmMez/IVmiLoYhIzDgob7iHAGghGP1p7e1O361iekQfBJItYPDnIBcCu5mTJ/uPgtefKl3Mm
KpTd+sDkTYaVAvlSQb78Z+iszs3/cZs3EgyuqUxOd91SRPeaVLXnBil+TMoyCUCp3CFlbeq1goXV
/79BAn0PqoZiUsMiC+Sr8lGkU2NQrojpxSSHp0gu8p5Kxb/2oLUmd+iTEPjU5Jm9QSMR7IEvetLW
ebSzfO+imY47tCC/TkzC4n2NI3JD0FwKUrEpG6sZuTFQhiCPxJA1+JJIE+mo0G8wZPUGJ51iSGcq
PmeKrg2lj9D5NAzFEMo/JK/Dpkm+PwJmnWn8kvHE50UBMflG4XkjAa4mVUy3wRDd//NAXP7yi5Ji
VLqzQKHrbqpeUXTUJ/nRKxQHL3prHBbEZD2C9rAtHfYCN/dWeS6b6HyYAgQuQE2QIHPWbhIHFJW6
Sk1THL+YQ9WFKKXJ+wc+y4WxYVn7NwshSF9PqcB+SlVhphTPlOFQojzN3aBLdA3QDUAQsSwmfS+W
Zzts42RCTqf+R6elYhZTkwwju9FbfdTAXaoM3d7yw5RHG1fPKYcZqK/54UQZ9f+EXJ6OENyEcPpJ
xz2uyGpKqd/6MklF37uV+9Ang5LtEufdydC4LcT5g7khHxJW108K4fA2Ax+EYoTCUiagQqiBjbqs
rBN9fWilvUAaG7T3ECInIals2A10xsiT+RqtCzXQAHLApyxFBvISg8BOOMO9WrodWW768x9rIjM2
MnTKX+KNM7U2jDe0i8qovQmv/K7z6j2y4EkCTm6zdN97f01oP7em2maVQhRsFSjEWk4iXP3p+2JD
idjksmOe7f+mHIFOpDiPTpq3/rhSl30IkHh83KNFtIYjLcOYopv7Bbn+xeqQPy9gv4/bNsb7zVYt
s//baAu1eGO3jHUVlgEwVft4xkesx/4AVd1WNuSatfcAdxi7fgeITNiMSQK5K93/DnJ49TJfbfbg
oddcCuWDlw2jPAExj61blSaxqx8Ze50PLg9b3iQ23YyNDC8Nw5zFULSjb2NX+6Giaygmdq74fAP+
8uznnUELssVYOWO6tyDTPk0VDi/ds6iUySe2J0ardCZKb6D92olma3nkhIqnHz+1liKsquapFInr
TTYeYFc6Ulg4mSb0dAKIYQpKq/D4bhkFRddEV8jkrC7tfhV0JprkdXEHuF96EPO2Doayd/wU2ues
gUHqn/SIV6r0QfaCJI4cXu/hHzMqPz2E9f54QPQTA0eC6xHC73txKPTs/VYYUuG+unF/c0gm9VHX
ljirRV3WQWqSSFr/l9R87v6wiZjxUmmn0V7hjCDWHONAD5Tq/pEjmInqnDUGd4z4BHjt0SNgCyR9
cLNegTxFdezwqbFuyp+k8puxNUYdvKsi4hbRwpNXCyjzOg9VTz+Il7WrF20SxNlAo0M5yVRgcl4C
VDGhkgx338voCelapx4XpyGVJKOwz170GHCNboCdFoyXSq02kIaGxUw2vc8OdCG4bdpPTTq/vvC5
AqxsZxXj7OAimjzYarznX0ppDvR72TbEUusdxuaEvY5z0hljHuSpvRc1mj/aPFFJe7hlAhWfGQtE
RCYBIljDE0d3uc7BRUMvPBv+h+85SUJiSTra3UhQR6Ld7hciqLJbWA7w+uGkikYToFJPegcS2QLD
cqCjmRC6vSNdLCtpWY4jCGQPQQ1F00nGaCzC1zFNVthdqJdGjDhnM4PsqfXiBi/PG2AXQ+UfZlpU
6B+mVxl97GMq16fq6NF40/Lw2d/rUr+8LBoTUY18d+IalGO8njjuW2ccHpDjxJ96W44Y+V+yUaKr
sAzJ1mtvxUHRet9eZmJulMD7WVCfdw5WOZnL5BAqyMxtB4s/HTj7ND19jV2w391FbR6s6c5iUmo4
vfvn3IDyGHVgqwSrIESBoLyD9VGd/tak7xe+MBUcK/HK4s/Owk9HPiziCJl/b7LDsD6Ygt51PL9Y
nX/MJToa1ufQW08qjpXCQ2joAMa1h6IPBUT+0ePbfqUQkwAoAkM2EBXTdkEmPXbvO+ArskWDPcxw
PoGx2CdxcRQb5DFdk0TljMLONm56prJScSCff7TyK7H1Ukwdzhc/sKXAaofj98EV2HdUFI7DlWZD
Jx9qOnVF+egd1fnO1HDdBa0e3rvblERsXXGTSLp2ekpKZ6Wa+3iwOkMst3vGft50ooYrGKgT0NHr
6e/g2TtAULGDFcTyaJypuhmnpWF3TPuhiFEQk/pGSnbVbHGCVDaU2TXI7BoVcgUgXaJZeadMJ2fF
iSWZKh7+dgj11M1nA+N6IfJfMHv4h0tYBLl71+4KnCYprq2t5MyjRqO2HB+Ze6WVibDOE6VeP9KU
bIqRQF+BPZA1yqX+a6KGDIej/Tc8MkeictfmsnvkALMqcAg08v5o4fG6KiKZ2ISeN+J4S4DYCq4Y
NTQEEJwmuTmgnQlj5TKFOM0saIg79/2FhZe3trU2Y/c9JbvW5jzLPPTACDfgsn5NAxu3lseNulJt
YwxV/h1AJWQhmS/s4hW2u4g63x+726VQa85JAd4HIO1wspQG3kFPOcrs3L6uGlSXrojOr6KzWuhI
lhVCcu2z+uzBvlSomHqSCWn89qIjBAdyGOLt1hd8GY5uup5vByAlJxLpKIK72ynCkwqAx0XH1byj
CLNzj7EMf16fifZejDSHPmK9JAEkqWH749msUCXjsiI8Bty55QCJjQZGQEr1ya4qfOTYcjuHet21
pcMhws9+PTqPN4mQUsslKlEz32+PZA0uRxpI3OaR6t8TKO7nmz5vK2z4NtbagJ4feg0Sz3CXS31E
j6Cdo+clURQjHYmL8WYgyczFEn9GOpVQuwD7IC+AwYd/TN3CoKTz5HIVmlTj0wM3c3JYQc1bxOo9
sJaxVznbDGvIkYYv2oBAnzLkMTuQ3uXoRASvq9l+VCBd3SWNzKmZqim083HIPFseb5uEc/NgDqN7
9evd6GXsTuTp4Alv/c5O5LYdpGUgLpK3W2aXLV3WKwGKAwvM2RRpEmqj20vHBhBg+llpm6Lo6y5y
IXqkrrpoNEVTB9sfy051LOBXYf2tmusg9uFguEpu2sch2b1n2uqCnEEDtxqlhxky609YkC83z0Eg
JUe/3ElIfZD1haxdhuAzMXVxVni339PDhbdiG3q/I1pgiDRC9oiyJsMKdVLWUykxFFd7izWo9aH2
0gPGawEV5Ace1cljzQ7FStFY93UHzU5ZKOGv2x98Nv7E7XHj80xwUrpgD91R4IJ6l+yLLTvT5bN5
G3bR35FPxFyUhnuzZpFOOa0KJJ6CyIsSZBOI+FO8EndQESvtmCpclVn932gUJbpuAjE5h1Vo8S4H
JPz2l8qtz9PpSvarfekDzSSBROx9/aDF+0WpverfYIyE4PdCuo5Hd48mXkbDHFM3r0qhzpF+b+AB
9j68tauDroed9ISSRLS3KaoqFvxBe0DyQfYjonGIadY7GgbnG5BBn4OPkY2+kzFfu/iRbHI02qA3
fve+89XNS//JUO/W5djb9DqsBu8GwTxXfCJCs8lMhDRpKZBsbwf7WNoOOvE1jSNvyc7HuG+a6tfD
j0bPvnlPik2nueMRB4BBeBT+NTRqsMh2K5B/JyxA5E8ws8Kuf+f4ylQcqgQKDAgR9qzERMAFwrAK
V3jfpXj8/JaaKtmfCEAqjgBHyP99UjWJiyidu1O2bxi6h+BXhnDeyKueUgYQOyr3jDSi0CT76ahI
SIs26LieMb7RJbdquyMlikKK52GIbYKATX4s66fUGopQbXfcelANZeeuVYHJNHiiwLQPIoLURVwR
IEIorWh41iVVz0Sih1p+2FQWZ6YHZm3UQBbzDCj1Qjz7B6xj6+0wF7N9esshU+rdA47afIUM/oC4
40TftFPb8HfG6ND9KFsygX9184Tx4/5PqWLRSeCdCljx/ag/sFTt0jZwF9IzItWaXX3kGjZfLABM
hiF58VHc+NdzKhoLO7y3TNY7OhWq2Ddr/HGplnSlSTQxxvMDY/rlyrewWXIPooyghkZ4gcCpIPEU
CzEuP5rTe+hnkyT3mnR4c1xVJGYQD89xyzDEOQ6ruQVTVpCxZPy7z/02AOG/YbRoifdyS4zLASzs
21rH2aNn8ZYnseaU3nIWI/cnRMdT/x6EyAJRpwshY80XBbuNfpi4RfDJZxu7/Knsq+ctq0+f7fgN
75bupW5T6k8+fuK8aWdo7KpL2VJvhtZOC2Ek/NDl3BlYLEbaj9pi6OzNXRJpDWJ+UwT4nJZCiGlw
TTxL9VRsx+3Ky1IylXke7drqFPHywu7WYfkvb6hZtIGhPW22WOePcbVbqMxeQX56siMBSuzpVQqk
gCTU8fiIjW3pBIixDXvFw0/mVEMS02FPkm9PuEaEaKPMx10a7HZ1w9/gaVFvgMHfIj8OhEVDlNdr
nUqdG6ClX3Mq8sKI84AIAxdq0sgVOZsd13elSRGdtVLWrREES8p5qV3S50GqOVpj3QTlAhRjV3vt
hIUtKKjgK64AcsFr1yBl3QRV8H9zY2uEPYmuDmqruForlZlwQmL4/drMBWBpozZTtGd0rHBZ4kCw
ogcZuy6kYFNW7wj7T34bYxOv9IRowFvGssHAobjKU4VqxuwMugCRFX21wV1+5xuyd+2N42QCUHMO
owqwxUxANSylFPdDcnRJ9qgES69Q8gMirjOATi4aObi+BI5YC0+M9gnn9DMcgBCacLF6N2KdVmdI
z99ISNwa7f9hjOgjzoC31keKzd4ATSdbn/FOpdy5d5hYiG/NoKKD7rZTED9z3jFbRskrz8hw0+Wr
gyNdKPrF1BkbEgakokbZWxSYmH1kFECVnCyngf7mEVqNfMQ7H1Z/yViJBdrEukwTUICxhRPcWIXC
g21B22rnK+rvRUcPNVK7p410Aol73jINm0usPn6ha6ZJ0TmwX44bQpTSQbleDKAwy7PxqjSVXW2o
6j7nIbHdnlT6joF4FZ+UZR6fGUg6swJUwcTupQ5aAXJP0FAeDBPuYlO/BjH6vkJjhDoSeTUv3ZB9
H4d5fQoWs+EB3vZ2HU/RZ3ZUOCXZ3qxmAPS7NSWNyedoarvLdiXf5kKPxUNUcLzTZR27FOEnnJ9j
KP7/M+EN8qipmIx9DkE1uj7aZYs+mpb7uTu7HlAWmAWv7UAuQ02c/aOQe6cB1SGVPhV7gY4A7qf9
MdXciCK+OSfeqGWOtyap6BlyvFZxHHbWmIpaK5amz3HTe2+fjHLtFCjk7ynzxaBgecF/T29yoVid
OZu1FJ7YoOmkAx6yyusr7PorOB05aB2UxY34bh2YQ/bukSUisqeEOB+Dni1F61k+siUJF8bPGEmb
ov2/U2JCeldLj7ZhrSbpjlUx2xjghTrs2UJbtD8cF+s7W7oBm7iePW979ajIVD0T4b0IuQTq5NTZ
gv7x5PQbnfnxyoBEnAVCDOl3Nczo/RLJCY9etM/qiqAOzMJQ1RH4Ze5Gbu/eKViRq6H93S4S9e6N
OlFxBW1Gk2L781zS0sSM9p8ldmh0PQHcegQgPdK5m5UqyFMNtd1V8WEVprN1RgkVljaLhnKbp+AH
dszjOtD7DpJSbFlTF0ihm/qMDkyutHr0ngVgACxK6AWlQZjaMQU3gggNBlNQVPaUjAtec5CSuZd0
jUEf/ocWu8q5nmgnYe4XaW3mFXrNYT+XqB/dlZ9Q4DK5KRBWc6NUgBZwo5PJERWh5CS9OAW3Sk/z
cXySjyYyedX7hqjsqvBOHj2R6mULX9N0XVanlabg7Ux5QekuQpRU/xPHqZP61ZVt79dwZP+lH5xB
9zsTzo/F9b0/I2wtaEfPb78rCv1R39gwXyUgg9P6hWxvvwVEvhkzfC43Qn/mw4PTs2UOKgKfgaKM
Y6ZmlVtWcKeNdlOaNOzqmfLmhkvLq9KMPsdZef2Wxz6qIOkihMiO+P47EaLw/DGwKRQ0ntZoZshE
Lxti8Z+/qqx/HzyjsKd5C/1HLgwponZULaTk1pPDzfKiwSl5IUWQuD2y3/XHFL2KQFUQ8H7S6Xh2
ss+ALEvWxTVMfPZzLbxpAm38+rEwHshegf9uflnsx3QcQuDfSOwbWTWyzfmxdE7M//YuonmNLAbR
lmsUAs7JotLlBAoI3xWMK1mhzSCCs9nLABzkQAfCJkEGud5UbTKAGqNaCDanRgdxl9VWDD7fAUS3
mHfabcfG76/sRTKD4lsXry8g2PXakOraT814YHR4wMAqOWNiL+gwgxLjhws5mVdhAbVH7P6yJvJG
XQQxVYLqIrc6DH+jyLLP+jky3kJgRZFXMyJIrpAiOFzx2uggUuNGIyYrStKKewagszLPnygPhSut
FPA36pSaL++sRuz4h2ZQVwNADEV2zcBL3M24oLY/xap1rqWGG/lUVpCLS+qjvnVIsHFTXwtBVn/p
OXuwB1ecBEa7vBBCWW5Uzp99VI1gA3mbr71SVX34xIa2EZNw3fiBeEu4hOjVizZnDghHvbpTaoul
cH8UoRyBqmc6XkwZo11TMKGK4OxbfW2vGbXJ6lTvTQGHju3v/9QCn6/ga+JOoRKbktJjArsEzgw3
RALlMJF6ev/C5qnqL5q9NzSOuTXo0bOxCsxMlpF6oCN51puA6X/rzBkCZFrnCGClBaHIPVCWklYB
GEaOP8HN/S7LoHqQf0sQU34WlyMZL2pPIRtlIK5LDc66KAuMhuRxqYKHEPbYpxz2RdnDzzms3IJ2
A9ffpH32+QsYcrkkWu/D9n0VrjxKV7dXRGWZDb0LAFNPS+NODLJ7+OjlYXx6Yf77wWZmgkMcLlW9
xi0/GVp7uNVj3zckR+ZMkzXOc0t1e97A7YioTqMMKug3yL0oPYNFPDcCkD50K+h0UaOycRM7MW5E
kQXsVgg7UoZg6AanbldM/QAKbaWW5L+FlK1d3VIjtEWM9j/J+lqaYRapRFnC3sBArtI9vzi3rWr+
RxeT4TzlNEsyuy2vRxsD1qQkrJbAWtD+TNOy8IepVkdrHhgJxOgva6kEffAHSqi/v8eap8sksGuk
Cc5k/QNhV6de0ky50Lh2+Hfi0+Reszi8mcJnwxUyBP0jHTVk6g9e7Sz1dDJ6hana1tBopkJ0RL8K
Vv0Lxdo1E82EAQ5cH5IgIo1DGKVxkrrqL+T6aLFmQCDxWc0hbjmTrNfqwlZZ4AnOS7F73R8RNmHu
8lagEqXYNjPth4AevCAbKcqiMbvRuZHYFCU+Spjpk4gOOS8WX/DfqGCAhqOQVNyUYnwDzZwMB8Wf
f1y9EsSEZVVthzz0ZRIsJfMlgrBbTJzD5QVRjPlLa4X7ACJTKUbDDa16a0cDSWpWWR7VqSRVSgVt
YMyHTsBXALluRWW52OCGzMedHqfrjQJQjsCOUVzGhiT7m04EAs1F5OFsshk5i5027vyvgJBiOPpG
r5Z++Yt+xkd2Ly9jQyq5gp6X9Zsux3u3OyQ1TMn9GEzL5iRoPtjHu56PFLxiNPRYxFExTsOjxaJR
qzAqIKA+LWHcRsMOiSocYCIgXw9n65q8WVfx700CRxxAXUaFCLW7ZNaQwfAVZjuj4sUkwiIH4kDW
yc4d0JbrPijUeBParY42iOCpkZt5Tk0WMHf4RcLMWbs4Tv36hMwL3ru7j4/CqNDa1tM8f4M4C9j2
oghdWGBQ+8lXI3yZWQzzCP+MC4LQekljhtI5TaMHQZveTDJWo/U7eZ8ZxLQfbtm1JEe59x20Enla
Flbl8k3F4jIeM655MOCNe8l8tw8QtM5ivSOkarQaaHkK72lFeZHExXPNbs6w17CZiPMk0N4aJWEp
Ckhpcmp2WH2JDYwNt+UM/eghWgwDLe4D0vYIOPXeP84LHy4VnL0sa/mREAjikBF0kUTj64AlkCpz
OOl5x2a+qSZ3YcznKz47uaAXpUHAW1Upg1MJb7vkK41LAP7OQdvob31KfSjDDH3BspI9kurK21Pk
CfNLh34Ra+WEW0dG3Pu5jGhgQnpeb/tNEQZKn1Z4uFrZcjGo+DWMEjkDo74JVdvFAY47WHuh+8i8
FtokXmBPeEMq/dBPv8Mnu3j2UHUFTv4cEL8Lda7chFZYHLbi9EcRjkqelHiQgrAFfFzlEqhDvnRL
V62ie1VptbtZfRmvtqRJhKwqH8rQpifU0w7TeUNGr5roTTjCXnjv4ap9Wz+53dJ6PX5uJttBj4jf
frg7/etNHLRNa3gfqkBp0hPM3BWtRcJXWs4KpTe2++yIQqw5jRo2PJx82fCcsJZM/KzRW3owRVI6
ngl25VIQZq7EhQOxINGizxzYQ6JSfOl6HJuVzaER6v0zNDpKXnicyquGmi/H0verGftxNprPyQ74
EDQxZPov0ILVUKVzufi+sUPOVUFHBCQVryNHsN7QVwSSlOQDP4H06rSF7UXuRPIiOIeWDQC7UD3F
vBgKEfeoiBSzX5/vCrcIcqP7BF2FAln+NeD4Am+FcWphGukh1pVy9g/kJw3OLlXTuh4nLONhBGuO
j5+p+V9GMwYX+l/dGHkT+pROWgIyj6wqyO2TserNu0csAyKd1p/eyk5OCcybt8VU0fXoYRs61C9y
+l7NOKyB/NA9X4fFP+NfqpALAgYFptw0HMZkvuwcm1gDq0kQEGFfLfjbF/2a4dU+SCD03GT58xBU
Ik6xI+5Kq1YaWavxGBP++6vk1PYGfgeBAymUvF+gD2kx5YnaviNM8VlrRaPHe4jBpIicmktjjqJK
/aKdOi053btScPmjYpPWDe0hV/KH7mrGI/viH7U5WpX193XcxDEpg2rYd7eYyhQ0p+jEvdV+Up64
dHHzUweLHWAc4nKSHFQXfZT6UK2dJcZ54J6XSireTrOHeML4LAQJXakxLVZ/U1togcH0G7AcW+9Q
nmAe81zZk/2bMnAiaJOG3BXL1hZSPn7LXf7D744sEUb6IFaYwtksjCZEoqeqM6Mb7bmD5Qn8FM+M
aYS4y+W9weyi/0G1kuJx7otgFUi8sMgclM1NJyAs8CsHqtwc7Ot6e7mrJ3oJQDuDTMURUyD4vy/B
nwED41xcpOMpiIphSOhcySt28jTRf6p7Ht0euRfpjVYIIiLja78KlFU9IwgovD6pqVVR1Ur4cm7f
gJXtyUgSAwcoqeSoAHS4/AKurATkDUaCBgXkBT29GWJTWo+Z9Oi0+YyUV+5gmPe62gG1KWZ6v+F/
QKGgom+36G+YZDGxKgSghEPqpqJ1B5khgdhf1SSJH9m5os3qvaMyKQnnE71A5unD+r41T24ar5q3
eF1ge9aTpj+Rk+mzw3P4ScFUQbw/ZKaM7scpaUP0lffuVEdJDx0Pl3ycB8ryNrzE1ik4ZJmwn93Q
wrn3AtvfNB6P/JnlrqCHZ9hGux8jxo+5fsLdhocBu9A3i6++KP40UQlw3j4/Big7hdLxoRkLxEpw
5jZT66IrtwIYmBF3Fk7nX85INMr0fzMgLwOjQTKB4+l9/q8v8utmOWSEo3SL0NVde0Y9xS5b3dEQ
SPDp9vkEynT1niiKBZBQshz8c4dI/eU4yk+oVrX2e8OlAZEZRQQfLw5RAPaXBg+0REPQph/Ojkiy
WOOcgxvQ4kUBL224W8QHLaSX36T2Hpmfn2XzFRsd1qprI8q+iyGBjNo2lsz12R1NHwpQdraEOE+O
yRfiJMWeMI+jzq4pkuuZJSgZMiUV5KiO5Nqqej3muaittdxkBbL+kFvRvxC3vMuVQfP+pePDJFdq
y1XDjQDcG7LPeK8XAkNoROEhtZXh2/5vdN5Jy6ywhI6MfNMPibFcOHZOaf7ym1ozJm5DBmV19NKU
0qvZljVVm5OzvbhdxPIJUa3j4RYgc6+W1Pp2BvJU26c9CiyXZC30f0WWXq+CCzoLeIyK24EtQrOO
23jnKwDFdpSqHEL4nlFvSV5bvJY3CcZUw2g4lHTOyMQVHZLpw81IO/Z0J9YMIMwOE+yX8q8qY+85
0K1WcLB261pjNN9SuiQP5kyjIai3HmdYk+GwTt6EbYd3/dShcIZEKQgVqR4qYXONAOS3gY3ras3d
ucyzr/YYMn8hKedzhuJjb/eJzhKi59Ar0SXeRclttE+go+zAFB45C9rrIlqsNSwJ5cj1iyRxny/0
5SKAAiJ1gkUuns3iBvqOYYc6KsZnitWTDYPEPQGIOj/RK6sce6Rkc6Tb6wqVmM1nxSUdhBzDU/Sy
Ayq40mk4gBXK9Zkg/gT4zzpxEW2EBxDXt5c4ErWCgdfPwiY0UkoGOlL7pugxt1RWRiUsb6YKroGy
IQMFt+2MrLSvsRFHgdHlIaxvfzAitK9C4JQwydd8hAsmRv/vdIl6b3xWH5ebTezrvRxyo1kTAbhJ
vfn4MwmNmXlqBvxiMm4auE2+8m+QWvABNuWmcPFL+wkWTQgFEsLuXewjYlaLxyPhvCCWYm0wySOl
Rxj0tJRNUYxDVP3yh2UaDyTrNqMOgI3rysSk/07jrGg7PkY62yO99smRwiHTAY7XEsBdHjPLWfqm
q5PqOD7LlWhe4vBZfLB8o+OxRk5HRh/dRUV/KKW0RpqCPoFt/OQ8YCbSjPx26sQ7FdaYJc7nWkXj
WyTe76CEdap9doM1AlVLKzdyRg91VqjlN3of85U2Y7gpFEEPrL5uwIdJCd1fL7sNiWSzLuWKC8zG
y9aXKCMKYPoIAZix4NocmAnY/O7LKq8YmNbME5xnZgBRdVB+YLxImVpPymQgEBJkpaq/HGe+TI1f
ua06TvJkvhtG15TTFNffex31Rt2cEVxVfH4dCbiTCT4X/HolXCjOdSAnMLFPDqFw+n2wkeYTnQB1
9vJP3oFXp4MOML/5IBFyfJlj7jqk74NNbtGAy/eKzm9ShypPc0fVIwZp+q99sZfs46j3TPeEX/9v
IsLxAGbDXqrVzzj4EHDF+pj6UZdvwUbDC2uGi0p/jj1D99bJv9R6WEH02O7Zj+cBYUre8koTL7gF
I8esCKHkfuPPJfRRPcOC0M5ylBNAEJv7J2yoNUFWtUem00RVDO4AYK7+AqU2MqEx02dv8elu3tv+
C4R4TmwTSjdFXngo+hHTROF+SVe6/Nz6UDryalSTgo32OyGJNApKVq34CiCGwUwhwEfuhOnfdQFG
g5If0KZ1Jh4o84dv+bBtHpW0timz49SwUDSpvCUECZWkU6MOi/OzLnY5lTY8mvlbAenXYicp4dqv
ermKs5AgqzwrtaT/GYj7yUgTnw8sa8ac/eKwNk9vQLIc3bwXRxOvESO0Sv/btr55XDhvXG+lJEaE
dJQi92qdH2omw5Jd3hk9OvwTKIcQlCdI5mdEM9HnKZQ2b6ZseQafkeu/8bVuPzlp8UXFunVMTt7d
1da0mWpvH/V8F0RVg0DXbN0WC9RXjGpWitsux+uS6JUU6eZMWjNCdIib2YozTmR0yeBYKc1LwmqG
W4MFzaz1adBaSslc2Gj4sADeVwdjKbqPGldrHvS5jml1pjUu38nNYZM91hA0O9WFaA4Ps/4pPOua
bppVzAqhOW02dj3JVFWxWHLeVrj7pRgr9r1JM01o8q8sNWlmhxKHcaHal6ukoyu7HOooO1r9R6bz
XxEH89Zu8L3z3EnI4qQSPBnj5coy/Ntk9NhxNY+XxEFe+0CY+vQ2h4dDsCMR1iObSXJjnvzae3VT
ZqTcc8N7M5UlWZH7um//tCaK+NcopSTXNvAYMsxBV+IZf+0hn5ghJirydMUl9rsMtiXUVEfHWM+U
nfvZWPqZnbe+XQUo01S1GQrjGipF3XkdJhQCs0+VPK81d9OjmgbgQeoXr6QQIes07Zukgt+nbkBF
Ei718gKRHnZDDQ/6R8Q4DwyGXEjXC8DxFEry6t/NGBlcnfqkeSq9Mqacjbvq378XjefFxhNGeZxO
A1Ae1Yh+xTP6Hzqx2qhuTNhY9K2ps7Aq7uzYMTRVJUHmewlgCZpRKvyv13nPWTL/g53BJvtoHlnf
zWkjeiHkOgeb70jkSXtvtTHLcAOYC50gXQ7Z4i0iZ5N9dE1mmKBjRUfeBYG5hlE9C/5zdnnDayR5
qGpt4PS2+C5yPuoNG/4CGdJ0Eul4xT6ytUOG68H9dXzX9rIOup77vc/jn5EZf/gtLuqK0fi1I35j
EGPr/xuHqhVlUsLA9APHyutrLt3rsAnvj8qswE2phPsIzDm7WYwvS8RyN9kugk62yEo4Z3vgP/jS
MUtHJ46NazWGZs1En7DSqzNj0ZZw5YZdiv/kaYDgHuXiqTKW5rrkOkmQIX9aiBrwhBf50FeRtOSZ
Jl/WVU/73X/rrzWnt95i0OzCdYH+CNBmg5nhjKvhsX9hnoHHLDYyhZ/dfMpMgQ8P44BbOe8ZjYu8
LVkBH4aKjqt9dYzm3jq6rA9GzOvnYwkFONX+wOAq2Q9QAxsDtnScVXHKOXcB8qov5sG8EWV6NnK8
ye335eH3nj0yi9LJkoa13r43gGatct4KiV8vY/iGRriCQmPNGzFpFbQZnJoLw9b4ark8qYJH+U7N
l6+KBNR5EgzGYB+4766iEEThyD5xc9UZMpoqdKJGgK203IUkKBD9gFhIVTNhoiiRQ1EXQBG5wiRH
1PrKl+bdIKKEGA9YdNrr4U2/odkEm7M7GlheOJT1FnqF4oWDlv9wwqYi3NYWsIK5uAObWFgh6rQy
76Ex/jUBqyx5lYqTRUjDR+7k3/cRZxwZAlFacPs8yyemWWYeLvMDESSyUlQye1pD5du1NIdA7H8H
ZSnnaxTty5SxrSXqJ4H3WqvkcyJxO09TeZZWFW0C6JmunHpVbuBpGbBHWrwtunsmaqqbPK49FFbz
cxu/s9Fazr51lmwRAyduDFDbvvTxfH1hpoMKm6bbampGwQOL5eTKFpv5CYoS5/+4RPn8S6IV94ee
6m+i+plSfYcWEvNsWehahZS9799C80Ml1oQjzLm2Qc5PH6ZrSzaOyjFoxB9GMCfIfHENPj8I4luM
hGqkFBRTr0GZHY1Q9aliYeTgNicIKc+G3XqmBgzdpK5F0i/2feC/KukER8UleJA4HEoL2qjlDX9N
dc6ADz6PAbCqS8+IKsD/SgOnFbF0NTLfzqWW2ha82xBVPtsf9pLt/Lbw/TXAGn+trTmo7BxuP22D
RuP8UswRubupAYfHNxOEHBuAyO9lIUIP16RJk9B4Xn9GIZjs6Qm2A/jCWNujFy1ymNkgKYcEJRSN
vAOBLswuyn0TKcS862ecPu5CJZ0eZ3ICplw5ycyIITRSIt6IFKQgnF1PuYMMqx22yG85I4JV8pYm
pwXB8Z9CBr2yRFjL8dS86WBZl4ohhxPNNm9D1XnuCHWYluTFluwdBmjmjlz7u8QV0RsPdvYpRN54
nNWUq/IE9q8w4YhCXe3oJk2cKyqKWee1vgbPTMi1IrClXLa07Ee1F7TbeKNeP7+cokWAwpaMUA8f
TgrH2vF1swO/MVSFRoz60bKjdPL8qp4i2tjKOgm5LZv3gRiKAxyM5M7kmxG/u6AJFc+AeztmDODZ
Dh11oRdWFNI3nqUvKSxeP6UsOQQwI/+V3vTn9v054vimtY8nSBkKuv8oQcGoBiFYL8d4KDaxVe2s
3xgmdLX1qQjlcEY/bPyIcErGg+lttHQoUEMUceZQtjUtkWKRd07rgk3loV8LbSLD7jnOtpiXCDIH
Huudkg7jUFC3MuZkRTBYwK7mgkcmEl6iW74yi8jQIBfDLmnsI7W94k+Mfz8mkOdwZQSgXsydnUIE
Yr8ar/VV7WXhHKl+2m891195freRNvoe14XYycj09NUOWhUA6oDTMugAVt0WWTRj2bp5Z4WJXG5p
YU8XY5762CDVB+U8glOZxWgzAhYntzKPKdFVDRLJ4k3O7cBR9ecwkMOy0niOX/bFmecu+MH4ifRy
9tB0V4c256TJ4DTLm0voJeA2Lg0jVThRI6IrVGMprYslHrkWOpbmS8hYXV/Lw1+2QigIEdYRker+
VJZLytmsjoEtfy05l0bZVP+3B047BxyX5Ms+iP1EQ4rkYSaf+WC32rX+PdVhEizASPGKRsHh9g3I
CVrIwtMaoiaK3QhzvmjSJbyO/RrUMDb+/Wwjzl8rsuHtKY0WKozVy4JfKj4eZiOZbhA/I4E6Wf2A
5HSuGqfqrFPG3d3RiV6S6CIsqUzWC0ljzZTknuMUhlw7gFstR8+PxIUvw5RZe32ECfih7glakRVc
EzpcmZ6aeC6U834CluIKDr8PQdjzk/ks534BwCCTgNyz4jUMVQeKJhV0Gnv/PZnkMocNFnAKbHiH
S7b6+D+Ta8DcbQtpyOjlOfXyxqedAuOLIMPCbeQGq4rfbHeMdT7nqs1kwNolbCc6LU5M9jyqXx17
zwgdhGuFfcrhMC/eTsJtiSQJ62xJCXLpkErlCgQKtQai3qcIX8RcA3o3D2ION58TIzqipHxeA6k4
XAH9aJUXLJn3IfFj24sOawq4Y40LCAj5RWXMVSbFlJ62WqV3U0lhYy5SvL69X6ngVbAnn3ym/cyr
nWMVc4DbzKJQilDcpmhoLyI/zZrDaIfdAWs4Q21oqG5ucqU9dnjX28fhObLonksJof0hnNV2jGMU
wf3xboCqkK40wIit9q9VQTurH1ltV4QyXFPNlV0027ftIxSHDh8NIjB0L7rOtO8cR15MsiIiWr8Z
9wYWWwuE7bY8Kroa0AmzpGYjum8ZVfmwdIxryQRuM0oPfwQ3WQJf6qNQ+s4KA0vKA+zNACty2ffR
b5gj9GwsA3vOxGAjQJq4Gnld3doMoKj0NCyQu6kU6yK8WwqYy9GBj60ZXdmEsTI+g2IqNByfVt5o
TtjmsE1bqyPvimoPm6sASwYQiyWyX6+6v2Jpf9D81/Z9pLWsIySrgrS1mg8Kwcqd3tZyX7LssdIb
RirMfMFibzn146CP+VhB2OYX6CjpjIqwOGSMPGR0Oy2dgNydMegyYJ+MoxaIQkVr9vUQ1fRUR0vL
bWwg9QWcHnwcx72RQQlyJSdlcFivzWnobQa9smxnbFChkLf11UbmcAUuLovXCDx7+R4K4fGmCniQ
DxAyNiHSct7MlNu5q9r94O9aktZI5x9I59wCj9N1OQtcTQ+0RwhJZEYic66cVzgAyamoS6rRrTpW
vdW2gwyrRg2w68dm53cnn2+327ruyBuOphZO9iB/eT7kr+RdVmlWqXIB0pUK1++Q4fEsH9QLbBHd
es0UhCXgaU3+TOGRKci4rtaUVAAmb4AOosaOAafD/9id/iEy4Ci7aWophLuOAtn9Zv2QUC1UDknF
pNvBULDmp3FPfPUtGteyHC9ZdwdUJI2X6y2ql+WAHE4DE2p9Aty02Rp2Xk1qLIiJTGnuS07X2piN
+2b19s4nDWL5r2xITeEgcTPzsZx/lp5IyAVNGugznSNe0484/ExzedFoVPcrRykvh0MlyluWUNSy
44dL2R6B+zyzStNKpX44+hLDW7mNdvUfiTk6rOH1Vho2E80umGb0hBpg4PJYqekVwYpvx86Jxmq+
AlnJV49LAIadhUSLjEOGbnaKe7oQkMBtGu4WlCCQSVwpi6Rb2ttVLTIihSMc+UK0rQsJzmY77pxs
DDBrXTuGfBbob8RNpQEWm89sqCUoMwfbvydvdbGpRB1VE9B6ScUXhNpLA+X9DqKKEYM0/VLsWDz6
0STi3PwVQCaUw+F1H3A1QEC6U2dwRrbaUQG/2dHMKBNdCg1giiM9HH1V86KUtHvIlMvNq2717gh7
TExXD7jguLtbY/RL+IGQmfiG7yHrGmW0mu2s5V6UHSIAyYSvEiKiyqu/WON+cy5L5Vzn/WfF6PWp
H6wqu27qqo9CBrG9q81UTloEZ0XTAJQZhNYUx2re+KKx94N5eTWSCFZ5WmFT8oeSDuW5+H4JQ2EU
F2vemG0hCxAm+1fFy7gPjehRGWeMOmN35LVrYCHYuu/CWx8mhjjvDTbbkrMhNc5arB8sdRzb6nhk
r1pUPovtM6fgEUeJ2TH+ckLJZLHjvABGUc5vgK7U9p++EJb1Ps0mZT6HiPQBbYL7MOKrHtrDEWpt
usOpyG9Pvzyr1Up9/OV51n1xA/IrK7UED+uj7CGe2PVNbzj6rzWxN0dzykeQtbRQlPXNnLpS0XOF
5oGTSH7/BcnwA+UBvhm0FxLgTuLh5xtf6EzuyO8Yjg+uNDvoYw3z8eRDBBQZycJGCThX0FcAjlyV
JNJEqiRwbNqv+T+hqQWa+dFlEboOdaBJAMdMb9QewW5jaFpDWk7UtRUkcVWG8d2GpI94TDT8rj6o
JGlqFeRR1sRO7jRAuwPLKLjcg8w5uPYKMJX7IQ0MYJRm5BmHnc2Cor424/OJ3JnUcFiOTQcAv/Nw
Uo0JYk9bohTJYiNRtyCO+7dsjDJhX2S0rs0Gfiwue5U91UckUwWGs70uwL5KYBwt9Y7XG1vUNyx1
ToYyZkkrhaYy+/zn7ugdFgROhOkjlYg2X9AzrNAenMYOZQbBHDR6MctqQXxjM+E965J/dxvdIA7+
kfjG4x6WKi3089yEojGPuLXl8fbSwEvKqW6N1IeM26JkNXRYXk6whEUDZwAuVuLPudo1l/OH+6po
skVh+zlV+UG2L+rn6w5yMWtFbDqWlCTBAxlvpIFTYHF4td54zwXCRgNsteNLcBercp8KldbJhn7o
7DbZkYzFfUTFo/C0pjhdkzKSpuoxXZribZFqOkGDp+IXPzyzVnBAttAI4HIk5oK3dhCSi+f/R/nE
W7F1s8fQ0pv8uYMmKYmh/eMHezRMPDN2cS11dxFABgP1as7MAorXRTUjr92bvySDfusupxwaPx7G
tq0oyHe1bxMnmu4uCbu3EPqGXfMAPa2fGBAHwKjqPQOfkfMzdZ+gMNJ926YzuWe9krCCoZGTkiWs
tAfnracGvu5ZahrFbSLNEbu5GloBOUxm6EQoDqbpBPptgzk2u6Rz80lwbM18nx2QFXYEKfSN7/iu
/wa4t5iTCXTtHJQHZTvGus9UB3APZK6xbA9ZUtmmWQteoUqya1mm+N8aUgT00eqUP/2JZStAmmgY
2fLFTOp/krCTQpN3s/+CuSH1fSXS0crP6U8esG5Nu4Ygok9fs2jtF1WUqur+DI1oOMxVIuXdHSRP
JvdbQnNnr6SPdiBrPyk1WmjHidP8XV2Xs2huGSUgvAFUKwB5ccgC8UCCWEJzDsHdtvZZ3VqOHabJ
bge6MhN60Q7bJHvl5jVgJV3bYfpH9Lq1NgWcc2tLIbotedFf7gY0kUBWJV+2uh4szgsyixaYk6qh
iL7ISxSsGmErj0z2F6YtUAIKafwtm3kRg7MtKMrA/qJwdi1G9Z/l7dJCSAcywBNAXE3HWERzGmh5
rpA4gD7KxF0DGK4FeqjzDjqZQXhRoWoBZV8ApIxPquGPnTqxUq8ih1uLqdT80rSu4TttB3RuZvzu
sejOuSDD00sX0gE7lMtVJXK1633iaxNMbmds512qI1ZmcqFt9bLJ25dLIRr8jIukSO0aPykobnvB
w/ydY1feTlQQg7EOmwR8cC9RVRge2EXZUKbPP8m7630Jty79cWnQa3Via+rkl0APk+Sg7ARGleZk
UulnY+MVG3E+MgJXVa37mVudHRZNGCsUW9Ez3X/LgQnanrhSOOUt86mX0NGaJdkPRNa5i3iFgQJK
ypUfIfSCgjOVX56Ol+7VAZzlC0KU03Bb0If0LH1zAcvWB1hq9h00EETaoxMxwCUDS6/pcwxhTNBt
lhzQsTSBJVdgQwp53grxzHrKHyhi4DKHskAN/yVMNxZUZ1Beh7SfpHmpWdiQwg/2mCC2UGa73xNI
rvym6lRx8DE974y8ZWq4fz1NpstbZo9RZ9SmCsFnnS5CkYQa3gl4tymM6o6rvokrlGqnR1Uhk6go
m+B4tVh7LmcF64UNyWznRQWIHL3E++7oPxQBQBXr1lYaZKvWx6jvSS34Vj/zxS6zk5q/hNJPLt39
jQ7U0RRGNZIpxsulYbRyyZ0U5U248kCSbgIJ17G3tty+2zVzvxS2zKxF3lmXQXkpftAK004//x+D
e178TtLoeOuH8r7KgFM7uzhC4C5nStKAKmt2WLPTlzHjNF0kgoRC4AuslVx592wGAf6TbiE+lUKM
iGgRg3egPZaINPK4iTVtCx7z21m788W8u7E1SHDFW3lcwjkILcyh74Lqnho91tueD9XpcfBH4Pn7
SMs5EbSB0JeHW3cvXZQo6V4+f50D1Da/AULjodwx+hEW6G504xg1D/aPkvkWT6BYgbRMTDqItyJd
0P6vDF/WBNzb7x0MAdswQAVUgyzRm1sySLcImlsym8c6pNFXI8VhsKRD+v5jXKjb6zzKBh6o1oTm
gpu+ZU9rxERRmBCqGXunRzo/ACRHXF6uVLq+B8T2uz/HwDTwjvtWwGLCuWIJNFtDTBZx/X7cUdO2
6tNR9JjYRKzRlNrbC04DNCgxTks/VSYgK8PieuPts/bpGitQNEblVYiHIJ2fwGEAiSk6qaTEPEdo
sD8B0+OhCXeh/AmIa14Pcqslfzw52AQZB2vvJIiPxeegWrX9LrF2dxDT4joGOj/Nh9DucY4Pw2pl
DesflMyIGvD0pt+h11K3mNmuiAifUFOgp/bM29AGz//i1TkpsWSOBncXKyYThitHiT6y9sOeIAhd
zwvz0iyYOsJmd1m2VI37OMr4IoQMJUqa3fTdrtXUrjo3cA7ouI71sa/Y86ZW6cD4FZ070n0TTlO4
uBVMKGqLWqwGT7+HMuqtD52za9k3VH1lI401h5f4RlXpI1PQWrQV8OSmK4nuu+SFczfHchROSrMk
yQF5xrmGZaAuKvwg9FlhzIAhSJvW1lBN1bp7+yhZX3h9P3vMXCgqU5c5bQJgOK/28IVWTnIIHaWU
jxP1Rumh6dsGxmmV56XOW7/oeY46k+faVjXKVe+AwRTnJi22nr4kWo9LyG1PPqgQSC+MmW4/U4pT
eThTU15/YKNT/5nyfvqXzR/keJRkXZqMmpayiWeNi5UJ6058m2vOiShHKx0HUezdB5TajvS0uDl8
CuNK7+hrWTXiItmR3wSsH1t+G/RUzjtP2qvf38HdZ+/Hbj+tgIXP5+MRWOyyQpsUUh4mGwZYvRAt
uI71hMq1TUWzKHI367zq3RByd8Gn2vUTpPMx8/7wx2ipLd2CXT2LSQ//Sp3zscJ2rN7tcBsA/B/g
irmbUbS9VY7F83Tzto6hkUWeTNAvbKJiBfyAF7sRC5kz8pBy20NFaN5jonHuWMZe7Eq+9tFRhSF8
npi2K9SG5CUqbKy1/1t3T+q0lu7gZ3321oKmo9mxROE1iBmfBPt26sjxk57clai1tI4U3ZRR5nC4
jhU+3v/0+Z+KDpMmxJu5Ctjx9PwRldjSqf9Xgpp9QySRrXIJK+mcPNhIVNQCMF0ynMh3ZZ6Rreff
v3yEtMEkigDhvkEGhkOLwUoZMBa2xx7SAVhlgyq7ECFFTlz53qK9Waht7R3hgJrgQZEXZWFLClxM
48iMYXr/hH1lBGt5lLJzfGzPFYcO1RO9lKm/qu9e7CxuY1NM4J+Bd1IS2YLMOlXwR41NIHYaDN8C
4e+9gSF7+Nb/+9QM+enJjWkoAdh+N2Z34ICZM6iaYYuOe4JdcgXkroFaRPxmY8Ifkp7bYXMiqBIG
rOcPrasr7dj4rtIjIdoomMn0plze7s7EoSZMj+Bh7wfUVTHDgLsbXhyJXAjbKAptYYaik1Hat4C+
Iyr8PRp+cAsmBC1p36PeDIyuAt4M0yxxoi4AWbtGpsCfNWdVoPmcD3OXsN4m+Ha8YD8b5//Kg1sj
kuBWcxydgMK+oUjFsb9aTbsCWj4V36v2n/951RIi9vxk5vyYHGoiUnZ+j5CP3BeF5mIAKepZ4iR7
p9HvQPVFCOVfdQ9CqB/sBThECw3+SHxt4VrzlFIFz+KAOq7cSCO+gtMMKhNcdRK2Hrzhjp0ifsrr
/6aLkDEYrxqeS0B6v0iy4+0woOylv97AvbJOkqeHR/ePzxp7PGdT9AdH6b/2u6HnPCSYT6vwkPyK
bAI+KJnCCQo0EQLT7m1wpSshpj4NCL9Sj+JSKenWfBG1jGyIHvmENjj/1gydj1D4SHEVxYeMQqtu
/j7v2omtTg20k9hvj5IV/9/2OdjSODD7mkozm8BCzjNskfeKDUgvAlCceItLUbX9Z0zf2U9+KNID
1IPaqE++eQKIVIigO7cZQZZWX6e/JA7Q4GqNlcUQpbjOuUCA5eOMOlC+8MJj0ULk9E9v4DcJxNA1
WQ5GUd30QueHIerrz4loWR+XISehn0RIMt6tl70r2o8J25UJqysbdFS5jf0JJ1DcqbPPNkS8lSAh
SdAtRTIC5VWcv5lvDxz8V66tKrFY+ENTfYufWtE4XiPrmMOxncADj8wBqCoU8fCnLl22m/wTAtbA
kFzQeXOjC7o5VAqB3HSCrPZq+exPpy3kyvAHH66Qd87w+d4uOCzxWsgX2jkZ1YlpIR/GWzkeNJtN
lAJnanRCMNhkV/n/jYsxQG/LJaOrFIy8HSbJR76Ywxo1sMbr0f3fYrxk4j7Zl4PmVp0h0y9Qwn3f
aGD2YGhMoEjoFHnGjfgwWFO5dAvG7NG1PKqTEOKcP/sQ+lyleYNB5rriWQgDj/jLt6dBgIYA6uYj
e1UTkSa+omm8abYwhA/uNnZmi0jFXq7LMGsrercPwf3LWplMs0v96jpZdvboUDRn0ugQTuexj4WD
SmSHs5re/jd/6grO4sxDz9Ad2xt8kL3WUGnFAXGlS6eDP4rRjJstwTWWN43o8eri787q7ZvpZWBe
imj6T91lIXAShJYdH177L+vVHIQu1nv+ydRwiDyOoJ2XVlRa5MhTp0lcE23+OJ5icttjp2B9zUhs
pkESkNO2uikSX6LnfgFqSZqICqfbKZumvyIuO6Lb8Xc+315Z926L06sZORgpS975E3CBib08ROCY
bVur2EestsFN8/cEgRdOdCRwHGljXYKFt0ZDkPP5m+NynAMw2okKQp3Yp/fdK4z9llczHttact9Q
aSwV443KE0oCSruPzclTZ7tlBzmrYk3gqg//nwMHqVWAgLi+koWTZ25N1isv59jNcmRQmyAEwsj0
guuB6Ca/QhWQGR6gQ9qGvY9OihJ2w+ngOTstwetyt1Cj+UjvOtLg8ZbWzz7B4tWK9JzXMSCSUydX
B9h1IinSEFZ+OotWA6o0VWj1VX7DL8krfhc1gG0pwxxq0WIldd8xpVqfEpgyPby1KPg3o/eqcKOp
hfAnYv4UTf0IEtiXPHXBf33OM+jQYIDNnRgHusPjWnQlHiMSqwOll2NJXGo9G1VezgTzYP6BwyHV
3DJDKJwokExbnNshCsP9eVCSrNX52u0R+zkvJmws8fSH9ZakiTuNORIn45k9eAe/2+2dsmnMMFF2
H7UDTaRnMnjT5ktXXudCrK7bu4bvh1tuxeEA3ZVLOyO1UyMFmtme+RNYaBZDpGBGimbx5kND5iZz
PfLP6NzBvnarusjmgeJIQt2EbRKcveNNvX5iLJRmGjLmmyF93AgJl3Om2BAs/qdAcptNwyH5ufYb
/vxTS4vR2UjdLvYPgsSD7ugbqSvpxisZhN4C/DJbhQKCNg8TtVY3fG5SAdj6Y1aEtq4mX2ad5rMT
0EfzFIzfRNHttfL15xsFSfEYczSXp2o5gOHQ6+2fQTgkuuTzHa7CM42JyKCLNVDRayRm7s6gQeCN
AlQnO0ZML2Nq++7I/0tiYkkytAN14YlxgxKYkIsgFksLjUtrWMQm/3N+gOe+GL9RIpTD425+sT7c
kc5gQsf1HbUT129EJjlmtfR3trYtCMnXrFxzqzG/rSHWmpJPXi/9Dw1urRj/axyeOXiDDWs5HnHh
IyXcF0AIQEQTuqQJQC/+0oKRjFiLpSFltqfqVbHvZl5GsSPWSxipFagvaef9X5MMmS7I+1SS0Nnh
en63TYI4FeBbsCrYgsV4qrEajG+C2xGs7+wtTzUNogCwC3rPakY4uG2L7WD8Cd7TbXA/0J38/fxT
yNC47c2GOHoZkU5uzG6p7+Bb5529pqhFqPeGTneDD0qnmgCmf91JgOZ0bOeuGo/mlTnjfSJMJsJN
CwDpcMiHkhpv6CY9MQ+2QRiphCdfHDcvSegI77BPO4Dfwxa+tWXueVvRJfga+sequd1nSN+NteXz
T3Vf1oUDxaLJmduY6HLhwrg8dDNsoiVUEzATbzakqPluvvEaL98dt5q2R0MDT5I7JIi3jeECPxmg
jXKPWKpm2G8R1s1r1/fqnKzDBzw17CGf2W36Uy5XJJmElR7KvzLNIyHSiiWJ1wYhAsZdgQ5Neq2d
OMOfrP/pHI2Bmf5oyj1+/ovr+c1PFc2O85OwhaS4efUYA7F0FUBb9WfSdOO2hTDoNhq3Pk7NdXEh
uHwGmx6tLUpR6lyQF3NamVuN1GzQOnSxoiWBWOTGBVKjN/zINp3aQSkv8m3zHZr+bnZRHPcHdfF9
gKVjooqtKUJM1DtMCZH1sSW3UtlQSMg+OmYO91iP+AAgK5ul6+dUyheN//exEhlD+E6Qiq3nLdq+
XG5rlATTqfE7p9bMjyhiMFm7JUCAXhXOm2it3XAsx5PYwPSrLgWKbJYy9BplojARq1V+hzPQeOsH
JWGDwHQoc4c1KOLjkkdcAzi/pcmfwQDcLx0tWpl+eRAAG5Vm96Gc8SiLlmrGVutH883kQDEml5oE
PGQmPy4u14GeObF3cOhCJCuIAAfg8ibe8kWAYyHPaWtAEFzme1fRhn4CTsXyFlFHze8hTbrqJN2j
VSX/Y0WRnaVz/IQGoUZ6BiR+s6rL5OXcPIZh2bdzkHEPBcVF6aF6fQEmzSuMXx6c+f6xd0hgLTZr
h/AoU0cTD7dW/QUnP3vx5T3cpb8o4+u9NGKILrRJNwnXGWX8KVtAoaY0KSb7WzwD6L6rXpFoo9np
D+ZJfDxy+96oz/vomWCIuow0gLCrjodAo3oS7GNVDkKtw6kErfPQLdv8Wk1GiuRCR/CWYMItfj2l
tY5xdQgZW8/QAtA59IYIbic1GQZRhgfDAXt7WUx37r4CptvI1U09ZXCZps+Aa83sWQL+zV9dgkFj
foLm0jaFO3fg++M1dviJG5fhZWyfe5zPLtN6KxFgdclN9Yv2BcupP4Nb3aDKvPcj6Z3DeqUDTLEj
ocjfPUTgugQ8R/hIdZ7uAPtQdOFaO1pIBmiAjMKLZvDsgOQg5dUP/+6wnvgyrhLhLcT+YCvmtgFh
25BSKEFuRDpzonNaZw8481bznQuLk4iZKALq9zBm1YOOC44HjoyN5N4yn8AKxcgaZUmoF8HYN1QB
NPhOBz88h0anDuijB0EoqCxZcrMqTi3tXyoxM/JgjCA6uU4TtoXwmW6cMHqkeCzMKLj2K/U9AyzZ
UDJ+mUWakEKJG8B9ghJdk5EQdLqaghRbbJyuDQPJovNQJZRx7EoW3LjvnJW1nxCTCoD/7d0Usn2x
3YfHn/Hsx1/Nu8UvUFOX3dwbA/1Gmg9JZRA8EBz8+8nJ3tpmS9eSNug9hMbTlSkfXSAIX2gchn8Y
ofWj5oQK4nyktcPS+vsF8LWw3UCwL7SMluDGMoQagJLVQOEo8Ri4UMfzTEVFfKPdMriBca/m4D6j
ml8MSCpgfR/kK0vDVH1XzJcjdTA5JCjjyDFWzVD8i6PeR+0WdpvsqcMMqhh5D6amHXQVYypsY2d0
XQ+pq48Kub/LsakGCDiY1Gqb/Y3dknlMRdQfE4lDSpGmQtwDakQ0Af+AQuVguVVlr6m6QKttkjce
NDPeTnCfUwH5gKopWLStT5QVpPbQ1ZeRdNwIF72Szd1gKJphk8ovZa5goLTRZS+2FBYlqO+0/l/4
kkBaf2d15iQXHY3JUUzUQF/01WXiFNepVq4eNbm0c8F3XZsOyMqgu9k3AIpJYtGoOrQtHzE2RDSI
oeBBpAgRsU6WgMkwJ0oKMITNThUz0lDDknzpu0Pj6EsTVg129/UhqVrYpBbZG3jPv3FQYUHNKWFu
sYcBXuzyy2AGuu2YurS39FzP5pzUq3Gh06s7JvwCIBj05u6sqzm3BIBZq7oR+FrQX5428Jf58vmE
LVfomIlAfE3fTG8PsKLnf6hY0H7nKRvP2dyky2bbAE6kme6GgDDu6zIl62UxczfzmHqkbneptqTP
+qAzYGGEJ8ixHJthuxVd7QxyLxRVYQJWE+KJAYmZofHqcQbWS6PlYgUNuZLXBDB3Pxju33XoWUZo
EzvibqftqoUw082+7FkfgaqEYc0hkFVWaXXz3T0/8pc+L2AscmOjGA5oDuuPdjchwlTDr7Fajuot
FgLd8Rn3A9Ind/HzQGzAr82lq4TjAiZ0SZbLURbnBJln4w21bzOzV4kL7GshUBK3mPOV5jMgLhet
5egO9NNZRLqtX2ecP9B7pwSCv7og7zOvJxC6U2VUVovyiXwIPo+PRPZXNwc9ZtcSA3b+1r2WA9Xz
wLg/nyUPF2KBDQFtmKTSD+2AqErkJ0g5ALmM9bIv4AichFU4nngmWfZD1ZBfGnp+X71XEYZFVLaP
cyqKvZlycQZ5IoPpCt94c9ASfe5tDlVFcjOCBX8C1PHcRPs7mmKt06ku83viyOLq7SMF7zKqDr8E
b/KQ/QVelJt4T7bbAg+Yt5uiAXGeiLKXEXIabkdzdpvx04DR3Q2kNwa0Tfbqmu9IzWMrTqgB7lwd
hxa6Ef7fcAR7+F4IKFd4+WCbpxeR2RXtNFBukKjibcRaybSs3+EUJdUZLfP6lbdo6g2y0v2SNTW0
LEkVbTDqOInVyCWxYWnVi/Y2gsxTAICRLWXyRkoDEO+kx3tmpFaELRCAzeWRGrXl81pfhStN56eA
DzCRCgRYD845eH6U+3HVdXv2xFhwgiSh4yBRaUCf0IETXx6o+Qkaw4LjYV3SOeFiBIjRqBQRcrvx
07RJqftdUqbLsxkeLUXtv93Bm3wLaXS375+/YvZg5RPYQygtGWQzu9NCeQnHBXt1soGXAkHS03+E
gHj/JpoU4QfoZ7eedAwYIV15pSP4nQe02q7XoQXnSSOL2HCkhFFCPjtpWi7j2/e4RXID+tWlmabd
ifh40YneLjoNV4vyDmDl73KcaBNi073XBFaMhB0ye2U4YgyCzaPYsAjiYkaxKNAQciBFg4w3f0qh
Lec+rkw3x939Xup0vXzVZOG59ZAzDSYP+t5emBK4/IDVeN2TSn+LPqGAzax2Xes0yNJ9PEbNAq/B
BktpHmA9AZXiD26b4CKjY0dBpGcKVFvNxNA15Dro5bIgW/mcT3sS0j9VLEUazDSmdx6Ac90xlojg
jQUAk/kEDcJiLcA3afV5RTFuOVWUB5zHFk2yy/vnnwJTtfOxPRt0eXGGXydlW41oA8bo/V+d+maR
6cq7lG2Iqamg7r53ixFCIFzjscY+zQ2ZARYa9sw4sDGDQvNcvN8c4e68YRENc/o3koO6hrkrEpsw
hrlRwmNCHkdzrvJc2ElY005r3lh5fYPcgkEhP6dETrez54Yy8//gUnHbLngfFKhf9Eg/uz/++1wP
C6sWdEcnN4pY5AXG7oqMu8IC+RYmKTOTmsIL3ekpFSWk9eLGj2bHGwOWx5KfeHecAwzglNbKI6io
LnloXFsjYUcL9o1gy4fNWv8PyxIjC98Dd/jraczov9sWfUCUfnI7Tmfn6ExerObhvYkNp2DDL08d
tIxICWnMQyMDbfM1tmcWj0bnm9uF1vOlhVGBkTzw/VXYYgf8CPT2GSV6ycmqJY0S3/iNR0E9gjgn
4tMp0kt42qMJ+egk9yNhqENT3lHUfeEx7xrfYZQqCXM1J2noSvV7dvErhXhgqV59SuXWictlFcXk
2s2nK/JqyWOgv8OAmyMUSpjX4Jl8eY3KCU0mkEm8vgBQLzVLy1alX5LaLyBdaAwCNBRTpbJE43gn
bsd1anAadB/rAAM9WHbMhAmdqN4xkT/DOrLYBOs5DR6MmcXuQSEsyHSQJRzJ3enA1sFez4q8E66l
ln8YGCfoeMwLSGyPrk0Uo8PgfRp89Kw9wruv1SRLEc8bAZuQ6OYj8+YyW2MRqrYXCV6nNJEBNXPW
0Iogsz/cNcHE/SOnEDU4kCtBvwSHMACWYf86kDuLAHV9DRxvfFe0hatfziKAPTS2HJ+9qzfhluag
aYgjbx4USGMburgrgNwzTdteMg23r8k8zqOn1c/bGYcShX+Gp5EBmYgfKyeQtYbiVJ9UZNWLbt5P
nQ3RBMUKkSoCFlwseCJA+UTPQ43W+KnyARS+qLA7xJEhSI2KUKiIarmvaqG7LJuw6WOYFCpBwvfF
8qzpF8LZdRZWpmbcf1ZdyWa7nL8qOpvY6hZtz27jnjX6TgRu/xRAy4v4pvIKkzeRzGht+Q/xqs8K
GtISCAL4svqS7CZ9FfeaF8SMnVseShEUlimkhrjuaprZJ+PDDVuJ1u4+u/H4qOqMpmZ20Tz20Or4
oE3zYRXwJxq1j476XF3zfrW4rCJgllNxn39ATy/3DJML15bi4p4PMMIf6aR7a/ZD25A4ADc6p9NK
Lkwv1Jwkh23DDaChpymk9DDKvh+MYZiIdnGWsKNQaCmBisZDktDlZiob0kh0DgvUyTGUAjSMp9pe
B6LMMFNOARdQES3qz4WC0gk3Dtn6Ot7r1nFwsdVu3INYMbQiiuj0GGWvYcEG9ivJXWj+stLqueqS
PJDF8LopLAviv6UVKMLISICOyyaN/slqDrxzkzQiKs+Yb7zbDVYoC4NRt8zn+YBrIsdgW91EafSh
P+1S3m3HrYJZZfUxZgn8Dk2T9Bcn/2urhex1mFVqJkTWgDAGs6RyGTW6QWXPI2kCUhMh8l2hPA3v
eMhedLtVsvwzB9EI/P63uYhVAnJT3xOBh6a2UQyS7U7EgB0fPkZzfV6S6Omc3pUqvS/t0MErjyct
3VQYHIRi2dyqcZ9PDnHcYqFJdVyJCIzt9zsbRFNTmexoxm3fGqo4yuKOBnZ1+PeSmsKQFpRSBLCu
xafaQF0JlKRJye9oivJuiyLYI7zSEd4hyBie8gUMqzHsRW+lXLSbVQ9hk8jlv4bs0UrTUZJYKpYw
59vUiLIX0Z2p09zwUQRRR2JFXUjmSBAQtRk/raK83z9qU71WriofyfstaCE3hjALBYgm5TPB6I0m
YgM6MmJLtUaI1z8AK/phW3P6lkefl6xX/gP97GFBOCmcXcjGw2qiPEx0NdhIJJdHY5wLK+5cH3wZ
ow2smvh6Gam+QwXYorA5WGchcduVDxCxnG3elDI0tBfnUeMfcaeheMCfNxPt9Bz5+wA01BmfsWJB
TGnb2vU4mP7RENzMJ9755oGiyWsTrhEe9eRD5vEpvSYF9k1hlIkVBOm5cpmOBcIaxZxnfDeVY5AU
W4DSdYQMDcBZg/PWGZIog6RS3sK4PeABbas2ZUe7AKjjrO52QQqnexXU3SByMVzpjiKx3fOl7vQx
ugNSPN7Jcegxqu6X0nbKFt84PhV6tLywgcVjZYOLvftRk0PYaOjHoovqyfVxt6kHKUjGEm5eRgJd
ZJyFwvk7WdGGtXyT0Comq8Zoa8GBMVNKuhOKUiyyuS8n8hYbbE+jyz67srbIzO+ISTmerz7+Eim5
XstwZwGBroyMTbQNufT5yKSocTlFTYa3qMGrvzx1O3jt32Go2DspxxdYq5+QhPGgtdX+FUkBFJtl
iGIX97C2R4fIdDUGjMJWbbKmFL+G9GxfwYc3BfWMoJt4GvX0svYgkkAuIDmO2jvZONoQGk0LoWGl
sZHHOrh86v5XiEX8WejOzd022B3BEbNunutT4Ki2zD5IUELT6Ar83JchrinpBoba+ejoqV4FQ2xd
fTrTErNHZ2OzwBwzu3b7+DfA8VYuo4pTn2jD4clvrdSWnVIlpbXbgzW1n5Ru9cQ/2Hc8VAJMLqEr
w6/EadIq+Mrj2MLdiz8EQoEZPA0Mrfrb5Cw0TdGLhH0xxdd41LxDCVjS3dsxs2WsTCTwRJLpIcic
s56kIwCcB3prPJ2dK8kjOsaMG7ty0ekCtvRPQeFgr4F9nIqFtViQLjf3IwLn9eg2yv5ZnEo49ELA
LOSjON5n+BMQvsysUkoLExXY1STijPhSEi7g09ohaMKAOrGeTqpY+3xUluENwjshsbuIdkj/OQCw
TCQyeKX2uEcwIL1AALxfi3P6FSXlcMTYhMaDHbG0MIK044q3A88MVKkorhpIO7IHNtcwYkJ9cnas
IA5hq8uHsgm7JSLhek9k5BonL+WcYnsm3PLOUKC/8ftd/IfAxQ8ATMPKvr5qtRhTmbABXf62Iceq
T10ApG7a2LC5hIFmtGnZDwiqrexxtnUmsqrr3dRLj1PUrzmPH8KKXiTmpBL4+ayVh+ydYEA0R3tk
CU0qDjbSjrQ9iqFWVtTTcoEOVMa7+ueYb6MuJqN2TtybrsdBb6UNpwPT28HiKiV1N2BENK3Am8Vg
U4oPjV6soIkYREzwenMpxd82MMPkhehFpKWXyiuTXlaF/V24sSk++6erhd7sH7lomliGXyYAYyeV
6gCEeedxHdNtH+ptcmgYu4P4t787/0jAFnjvbcAv4C15luUlI/N1ahkzbelQChLekI/Hsf5cGK8o
rjSua8bFnz+5sfIjI2EpDYkoXW6zHUbEgsum0zsL7CnIW7dqqJLUJ5z319JMvGylIIhrXaXd9S1j
zZlYauAdUdVErKZwbENqEAwXlabM6defR9DGRFeul35oDCZV08POlPYcdQafjqoEP2AZYTITYYSH
OVa3C5m/m1R39e/5yfW/Ry0gY3+VHAnnTqaVRj6JI24LM74X/v7+OIPwX8j+XnRGqhjYg3rqNE/R
5vviKyx50QRozDKw54stnzn8WniVcw1Z/09ox2dszY++wzoXz3fHSeW5qapGesz8Q0Thu3DT4n5u
IfaGSCwd5+4YPBW0vuGTjJEB434he2mRoL50GjyTdbEIHvAOwqVvFSvZpp34KeGXQreErtu6egCj
kMsmkKKTRB0ptVdM4wYR7XYjVQWVzl/pemlOftx4JJcPP2KLGg6KVV8cpQkrL+mRXyeMqIk7xa53
/5qIUZ9ECs/G6MuFU8gUtW71gLhykhO3iq9tGNhU2I51pszGCK1e5yr8qthmqhGAcs05H1BBYvzm
991DRKmqgK/pyvgEQUJCUuZ1xuu9jmUQIslxtdIpJn5PkWay8mFcz1BSTVUnOmosWi1JtlIHUeNx
LwYxyhVsSGNFOI4pdu9EP9vMYyr0ASU3lsZ9Tfw1JCfJ8pFb5KFWquFerLWUjAkExO1hsvgL7CLD
gi5Q/S2gI7111GQKxgaoGPSNKW6pqu05xKnk0qjaS96QNZm3ujnGpwIO+yHElmVs6JAAKzOanjCw
7PVtY7WAYmcVAoiOmLattgrBl33UHJdVz1tjjlx3EkdQtuxbIPJBnMVZn85M5XadcOHrB/ImdEAm
R9gWFdpBIavI2uUc4gc+rdPPBdOzZDAq3POhGUocJGtsBs2r3LbvL6591Engi6pDFtAzMqniirXR
WNAFByD5AGUJvjyBlDKkZeFEiHP5bYG08c1VCClkBY7zM8AYyfTYAojun8SU8F/OwjM5g7ckp46f
6gR2aW/RZoOrur2b9lG0H+sRdXf82lEDzBAI9ZH+S1zb+CEaQGoeJzkPLXzS2NJDnciLFl5Bjqwl
TvnR9cWCV+RrHzrx3owvGMtOzU3RHqIYCfNbEqAP8tEE7Noqor2ZQUkJ6s3/lRq+cw01ovl76aUQ
ZBjWc8e1DmWUVgsbm+lJstjV7vh1zUUSSFQX/eVUETNpQI/UVVeQfjFXy/ICCql2Wu1fY8CZP9QR
eSZSnuy20PZM946YL2NerMld9Xs74i903I+P9+wcI8oupQwhC3u046/jZU5iJgYytEhEPq4ob2+l
HsNa+XfZdU+/cC0juEUMymy5lnwBD/tLVNlcBHkEoTaRHAAsL4sA901nu/sJhozgB57uYLujH/I3
BG+PJncSVOo1pppZjFitnnsXCzmUZARoHQifSW3EHu6dWfT1D5lYlC1QSoK2FxJhlQFz7hh/fAUc
4rzQkbIs0T9hKtnQqbfoQye5Dq8hTpMhDLsIuMJ/J9w72SP+Bke3vUFCGDV1evYgYkS2NS73jZRK
odvvNX9w8u7xn3nMgqgjDI0wT/oh7mXPHfJLt10+9556LdB/QLVVT4sp87kT7FqTZ49GQZa/E6ej
PXXxQjcOwAqaDp+vBFoXCUmpvDRFsmVpy/00DdGRhq0ABsaNSvLIr77X2wmBNuHSQD+SuPyi25BN
yVT7rnPlp2t+gTgzoik3E9YFbsU79kmV9c2dOmX4+gmP1d5Kwdi7syX2AsCLOJM8VMVnJ4A3PvNN
MNm+KnIt5dXgQUvlc52u8xV8yMzvEgKbCX33HZMVL2Hp6aoh//vV/1IQiyjhm6kq/ZTEqmtMVayB
r6HCRCxgdAndaOKic52grYSqkH+ZHwSq6Jnji0Lr/sFhn0qN1cL0pMdQrUISNwb763oHs7OMG5Hx
jNjHRJ1zLQSRf4W/Vmd7DNA+UwYtatYnUQN9zrgnQlc8+sKcbJHYwvyyYGygZNG9wcm0Vfm294FU
Uytcemy2oBGYvVwt3gTgXQivgMlUlaOdw18b3mVpwuK7a0/iZpUiYIibrQhNC/nrW/CSN9zU4kuE
bhjGl0eiCQT5bTGYy0LgixjVaoH2B/y6gjHv7KuJQ0oEmbw5RL1tMpRL/KDsjjuCLPyGHS2FQKKn
Sxa7zvjS2gYJrsTENRVsgER5De55+peocnVkWmrMQkZLDhqcmMRIKvZ0fMmBPiDFKHEmw4MaMZOR
zo73OvS2kOsqeZtd4pqPra+1xOXI6enOJaQtacSXlauEfZ+ZDpRtSEw7NGemqdm2R1S1J9ojqNi0
+k02WO3FaDwdybIMkkkK5NdB9Ot0ArpOw+XshvRz4Zo2PX9OTMJRDc+xQrH3qxb8d7GAxsKiay4R
Zsry69ajKe21e3yYly3KrBmkfcUS77h4RBsV5hWyx5D8U++kiDkmlCIkpMk2QrgeBz4YxWkP5yMG
sG47uPuNu39MPilHKamdl2NNQUkaLyc3ed4CYoEcWU/nn2XNU5o9/VP8y8M141QhFLXHqMxl8Jsb
rH/3A8ub2HufKWUxkHecINZFZcWXHBU37lOfw5qybRt2lHqkLfsSbdHAfVZ+G109jFo7jZc+HALC
jWVkErk504S2qd0m8rsSBLbaZphW3XaHjTIP+Y+b0PLESjGYyi5xw6YWR/qsQMdWFCi1/wbh8mtZ
wgPLdH4RO8uOXHoSBLrL6ZW5VlDsoZ+G+SbHAu8nF8nCJcaevA/SKSpBxUB2HaRF1FpKVRTaz08p
p5zuJa9SftAcp2Ym/f3WM70YLVIg68rpAXXeH3wfNr1eL1uHcw1ygNZk+Em7QLuFER3NkIys8nMm
CEAfAyo1Hwv9/0YAjyiPS6/fPKrIpgpfonEPWhwv4jXD7LP29nLeGxU65ppJU0kFfjNLmFqBqqbR
szCeyyFkEQHmCr1CzMTciCri2bE/UR619BLUK06PFJsLNY8rHzPUHyYPtgvximcNsZSDiFzr7DL2
gF//9DRmTvdxgdlXhF6lDVYXfTPh7W5GpYUdKwCS2Ipm5RxFoPxQD7c1fVuLDucUqB51tKpdX+pq
mHXzt7cKiUeQP9qGJ2QIB5PTSgLZTlxNnNRzK4TBqCNwgTfVkzX/1Vk8SYLdaYX+vq3IdV3A/Tk9
1wN1g1M2C3BfGTZBkmC3iuo1U9bDrS5EdBq7PZEth5qEty12oF8A/1c/cr2IE1/s/0WSjuESgB6n
N0hgWU9nRoxVFRX6w7JyJT8poI6fBl98ru7a5TCa09v6z3JXcRDSUMe2UjSRUbl6iuPbsKcKKl72
fP6+yBrcC/iwsnDJwDO+ICTQYK2uMiuwMuY12R6ASynACXde6dLW1tXNsjV79qYuS3vfZKeRO99Y
oJGzbyr3vDVR3dMOY71lRTXohlJW6GwN3bZ6TeBR6q+U9Po0kR9OR00XnT1h3jE+Qrudk7erh8lJ
cx+TCsWiQctbaYzkqMvqcQ6iMBQjmceWEkiO7WrfzJ8A0iNfgXjsU3SgMFO2Zx7u01XCqLsrYLGY
zN3ONzh3+trQ559W7XkOz17fi7uJJ37aHGKbEIEpi6MTpMp3Znxeroeewjq2nKnRj4MTZH/IQ95y
1JHmxYBcLr70Pgxa9ZtbQ62CmvUx3bkPejGn/hr3E7IJ02I4kx6JYeR2QJE5KRuKnQXx9LipBsNV
daeKz07lYAT3HDxUuMBVul0LsjSpz1ZMWnQxU54UgxuuWrRuGp+k6eGHeeYuMuWBQcFrJAL3MYve
340c6onID5up0F8+URCUYTPM59hGr3+s/foKeyRvmv2xcar6f9/no7odLsFpIHeVl4MxsO0LLV2z
lwW+J4PmDRCw0uct4/f2JFm0hTl5u0ywz0gkLUz2byMraRl8ZoYY9/9KCptWlrx7RFlwqevUXxxW
2JZ+9HPwlDDlr0vXjF9lVIf5Xvyo4ogHf/5bdQrFwRIfeRvb/W+Lk9ejHxaZhlyYFWui+pGrd6yt
MejeaBHubdQmS6PdjRvwK7a4YeQ2n0+704j1fQ/ypS5B5XKFrn229nQssGZxDf4U5zZY2CMqbUEu
jBejQD12FA3N/TJA5ilRVJFb/30g+157fWewO97Z5wI3ceF6P3uXIPVcQERTnXP7/DP4A8xkiKtF
86ydWLIhoFRYV2E/7Wa8ArHKIOfdR47Ypv3RCbdcXamXT6Wk6DO412p47I4a3rPdBNRrE70iJ2mW
HPROSwG382pu6cLMgDwmqdlYyhACogh5mAiG4gpMU1IjnIf8Vso5O+uYNCO5X6QMvUTiDmF2cxzO
dT3NG+Oqeqn2hnHOhhuUIJ9cMRAGdx8mQXd54lvUsPEMWqJb+48G8XSxmSH6xxDy0J8olkja76vi
ZGc44zYa4WKCnTJU31pBVKfcNyXeGEe8duvz4T3SAvu6CL3fo6OdZhht3IlVmcZvnihFgw8zVfAy
G3gcc6QWdMqCC+qm2iQA+M3v4B4gLGhxhtqiMzTNzupL4IWh5Y0hw2jLtkkoEc9qiBqgTS4fsQ4C
UUcsWKnCHhgl6FDKXQdMFJw+Qse8lXTe5bGqg+Y6TOCM6oxFSkX9Fgi0mUkMFEGKb1jR8dgNlQQ7
re5YLw6oshezPMVPWnHz0CBd8EPMO5ZlVyLKs9mlFe/zQl3ogVzFhi+K+aAz4d5XVmPdxm2YbxB9
UBy5dCplGmiEufPqBpbpbIk/HKLL0QR64GOfmL05uihRsLS5AU4dsvZDQgc/gQCRnmy8b4DhHNF5
kMsS48+L4YKeULCmVmJmMQZGR0jthw1ZsbjoaKmXkTShL75FnltieuJ/7JU/6uHXYOEQEBqhL8SM
e1uL/zJlmp1qV5ij+tgi60yF5lx+OZMnw/UtL7mDKa+aV8NO9tax8lT+ycZFLPKsLqTDbmHlqwJJ
7HkVhWrtSqamAOdpNvHI3P3Asa44DXnuJDDO3QvkK0qRQ3BMHZdOvn8GXS6vWnuNCx8LJJ8BEksu
pLL0OB9N3WS8ELdipizRY6nntshq88wXXvtnlgPMABPtVFnC5dBczDgBgTjuRBbDvqMWh8tSv2ts
eMVT15PVJqoqphS5ys62ktkhSvRhg8OCSSQ9j2Mgx8iwz4UEo8WC1El3tIPHs7NNn3wOabISwc6E
3Yp7LvmDRJ4ja5mJ7DMkNk8Usw2m31mL/gq3Cu9HQsN3hNyBzdxsXogcbVT0xIXJm8fIA+LBi3HD
sudR6fGLRYTSJ+7VB2v4YH+wy5sOL2AajJ1fZhzRrlsqaah3ziOa2nKZizDiLeXuqDTGuPXulkok
y7HR3E2xHzyX1oVSDhLSCnkqbirmH4MNX/KvMzCwRgkcP3lAAtmWm/zIVu27xAou1cDBNPwd/Kr0
Hd255pAsoFSbYFo7PMdgxDEbbSVvKPwYlyBMNV1+Ef16xH4JYoy/kD6emnJcEbbIsd6+NbR7fNRI
JHaRCJfSOEbET2Nk7cCoMKCYMhridff3omF6aCRKYeWOTA0AFYJE+hF5ura1Vo5dFz7N03J6Zqu7
OkUsAGlQRW1+P+Ad1f9g927DbFEpMegz3O18wjH5BWmAGNp2qY1lLGX2KY9SDPcGnBRhZFizK3i+
xSyLey8l+pVNtFxcHzN5mC54EyfU02iclXDJyQp0N0/hbiFwWol1qs37q/2i+XXbxNuobTRolMd/
uosJV31/ldB6j1nNK/7PyZUHB1WruMr5gR4E21z9yBldC5rAgY14LY2KNJgC1Nz0RZRNMhEOJ4zs
aFu2ib93ry4nkz96uTIjbqx7+/Cy1GMTxEf7G40v4F2CQXG3IHTBNB2McPArxLSzufV0RIOvV0Mz
T1sxH0WZNJ82QMIsyifFilchMT7DC8nT0kTJU3rGyx3BTR1UlKjibI+JytSH9k4l6cyobM/SnKUP
4PdyxcLwwf4+gkCIKSkzN3/flJ4MBL8gZBEPldBPlRmurUi5CcmpOkpLcODqBfxg87mKZPvwLYWD
v7pcdgb7YJYQ34DYppeU3JR8Q9UWOw7vvLsGjp3OATP0TS6KsvHim6yWKcN8RBz3ZybAaCduv+ts
TKgOS8dz8yebKXl6qfjRh3xLw4cAQuvo9xvw3m8aSCS/oWwiCpDE0VwmFcLPxbGmsblSSDFOUu4x
6TQpr4fPPAmUnDBu1gbAQvGwHQNfdhd43GUofZp4/3mWoIJrJuJMAb7mDwyszqdmbEOWOrGXZ9T0
N6ZH1yC8KOXf9B6/PKNDsYQ9C1Nr9kLRrjTyhEq2vyuq/5Bxl0QYjTiUQPoyKlfWlN/OUWvPZ5r1
CLiaKOvD4E8eiZUZ4WY4wfG2jqPULqBjQV7Q6KztzgrHk/0I41heUs8E1HjNVqRU+tfotEs4YMpr
t7SM4X3KJtjvYH53ABvf0pFuHCwWRbs6nVT5lNT++0NvSdwv6Ndrxku/udveUKlyRGTnps2M0VZJ
W+lA8de3PN4L1WNjX3gtGSst2qKPsLPK9SCsOwS5vrB6bS0wCI0to44Y6/AyqqkIAe0UVqHaPoCd
3Ob8UayUjSeua6R8OfDIHZAFjTPQaLGPVLU75DJ0STX8x4jRQ/23kxRIbcJ5a5lx0FUqzVapyeeL
q0pLtNNQYwO1LAbmrfRvWOZ6IIzbWZyCe/J+A+H8AxzDCiTGM5if10pyXAK7tkr9UHErewWhijTz
Q6NZYbAped+f/tfXS/ZAmVl1ABC6ecjbWYOdYMdzbIN6y6KETKlVGc+Nbh8GsQmYmajLBByxnsSY
5L9QWCOYk+ZQt/F96XlLZcowwRXKYXRBO6KBYVT8p5gtsN8reycj1GK4FX6XltUDVuY+L+WEq4ms
tevD3/2/StmPjXDGebW+8YWVbJvk9qwfnNzDzxkqigaYDLIpI8TzvIYl0wceelhBILl+q++R2GGG
rh+dvFFTjA3doG1L4Rpya/x8FTXcTPnWdFd9zNLz4DZFD3HW3AGvbTUFfXAQ6YJ/0lZWpKRNga5p
frl5i7xtLngMlUWpSz4KJwGqaWmy6/W5e4A/D3WVmYN5UJ6/mxh3swjoaayOcUC7NaAlvXxqx7Ei
f9qwXE+rLZgrXW3IzSR4L78obSY+5vXzXz5Eal7lqHiW5p3x6rN6XCQ8lAciT26d64SPk0KesNxq
Q92qDsGACrzooCAqjaiCu31g/e69QD/o6NgkfhPjWR8agX3P8hnRwBJblp6YqFW3SRroEK7XM3D7
7ZVQA/wpd0ob1tvKK72jLNWPc/7+Mi4h8OyV4UzkcBVuwxcCJRv9kz56aXfR1VxQxPx5ZAvJpLfp
PHU+vPQXGyHkdqf/MPWonKXaAetq6FUoULi/bIUuHar/Cptoq9KHstzxo+vLq7JLQ0PvFTPGudMC
2O6/PA7MlhIeHxhuyWn63rH1/JbH89gxFoYZYizjg+mXdt2B1Pe641dZxjRcOpGxnILIN4MHyhMc
lRrXyhVzMr1hyrH9oZiF07xp03cTy4Nq7ztpskn3/nay5e20QeQrNpUsq1g2Hbn/wi+/AhcRPabO
nq7ltv851x5Wngn4KOz9iT8C9wMUMNEOIWK9tLh//tudibUo1LeX1aBkguONyP05x1RWdMOwRsFd
rsjBVqcqreimY0uNK6JWFKfB//Xs/kYXnw5ttXSNJkGW7Bb75xmQIno6MITIVojD+Yt1AMIb0wIW
hXmcXP4LRymDrEb2sa2Xr/FbGbFx8Por4WRDYDXjFkWBIodilr6Nv0+iMRcBmHznGy3LrrHfFSZN
cydWcdXPSEQ1PHhQNHLcbUKymNIvREOYLnGCt75qPeV48QrVHL/Ty9udng8BkX1kkSL95zoxQSyE
24Oq/3eLiheFazFYSIU4/lk8i3VSL9pMTIxE9apJ9R3brA3rmOGWHk+p/ktOK6w1Y8vei/gg1h28
GlyUySJiXw1N1UGBBns+ssu7gQ7C7zbWnlmEBa3ekC/+xnaHTeWp/l49VPE2a8S0e7rTwtHSkQWU
TjuFiUa8MUsdKO7J93rItRiIxVUf4C5oNWfz9lOop82Q8JwdrYt9lbTipujTtxwq2xzzkToEwdGH
/tA+4l6K7UMf+JFBKGC8Z4ZatOYZ6HISo1hb2NdNAzwnxeoe6KATPkw8+sl2Xmwh6Qk+YAT6+lif
5/TwtiqZa23tQpak4VJxLInUkV8qMNEKpGV4Ks4vOSVXhUi3fOTM/fSyeD2Xv6p1S+D1DRkFG0oH
LVrveR1KBakXXYXhi6ZQZdhHwtPP1v9ExxZDfk3XbuRWfR0pXEk1of0RJJiz5mgc/KyzHIvMe6Fx
Sv5rqkb569NLMK7rSmPoVpN1pEFHaYhKCGNvvu0x3uREGneXCJ8bE63SlABWaGvjQ2Jhth6mTicS
tkJ7vMjS2tGH4CJ7NOWaYRQ7sYSv/cms4/tY2zlousHEo6h3ku8CQnyf47RXwnOXJVuOlDwUUea3
5gOSeKP0Joh3w4xpICN42Tl9M1lQWg6rTiIiMbRBJ8MYoWdUD6fUbkBj1RMg6mi99JDte+JrIBLO
v5HFtJBkuOQZxfrLOFYDEKTLdWnI0epylvRdxWNuzdtGrKoO7voidtCkBPeDHl0ZBnDSrNjaxLe1
kiQT1AmqPOVnYXDJ6zIAQ/xMaakiAqTeJhCxhl2NEI72h1AYbn1GfdNFK0fuBg9mW+on2i88C6Q2
2+zs3L5YDWHD0ecGj6+bqGzS5LEyumQ+RHPBm5fCUQ+AZyQCyLo4yr5hQLvsiecA6uXrlw6XwXAl
rfOTNMtVUnBRKnIk/XgERqlWwMXZZViDalLCWwueP8Uu0jYwez7IhkE/+50EayDasBM0cwRt6SF0
1aQA8sqCWb8kU7hUprFJD8DtCdbS+lLMvUdtZerR3IvPeWOW3Gwc4bEB3kIfCVMaBlmPUjCjrv/Z
ID/+HziSNmhp4kQgxLhjuSVW8g8dMJfISljH0WdSXiGTm7vfpiVs35nCrPZxJ+7ZhwbbsBTTuLLj
l1cZLyBzuMMEpLi9ox8OnyQMCXedux/S27E1hTKWpS0J5iBMH0TSKWfXlHk+rZM0c1eqQh3hP5UY
8EKkhfbK829Srf7Wr7INTVTRxBigDl9x0S43a7/lV8Qxl+Rv/2DWapOMIkN261GIVncbSW2l2Uyj
JYjdOyNiR5L8Cv/ex8S13JDajaTe0uPT9t+r1+GiPv4VnXE0ak14LsZ+uboX8kzv4o29p6MZUch7
01lOcGtzz86YtqT23n4cOG7hlUla5lNwR36J5f1asIV9WdmNSHkqPGtnNQgfcys0pxdZdGVFaf8e
OR1LGrQu3fGv8mqTIhKOnLaJmYssDhBFI/JUTol0mkieBypBGqt0J8zHVfx+/zsWDSyxawM3w17c
I88jwruixDr364T+34k3puzMNrShB/qDYJijKRe5oJQaLluzZJVjwqapHtw1sJBZWe4BX4Ccullf
NjXH2e/5KBiIBlU4CjaJ8+/DHrcmHRRCPjffZgjNtKuxKR0gHAoJrNFtnqz3J1KYuxrIBPimQjBF
hINAEWax6c6ArEF6TzPLXxkrHS1sU17H7ijgNCVsTe9SBaySg+OmtoEnBuYXrbv7ARo4PlQ9VHFb
MsMivRmYx7W9gcQsTvk7zFtuOBYPq/LT2eb2dcfgs1MBHyn7v+3p9VpUIAAdcfgx11EmLdIGQJBE
pLAwBtEhMnuZayfybdbkHfRGuqRXM+RHweyvX3cIsgJGOrh4RmjO8k2TkjgVK0EOwzH/S9IELdTv
OcceGfi777LuwXxchsysEq/gDB8xPFiUUf33OjnXkXAl9SMLKIyzXH225QcLoTEmc5Ndmp3WyWWQ
hCLnav2X2V0mNxLUlzdOfbx3ZNN9x1WVS4qm2+yARKaaemxWZWYQ/eGD4NLnhBMy7uurLEc35CPC
WoFv+4jHvZO2iPpPICF/ayEQhSdrAIZbnYov4iPhSzmYl+jo+Nps8ThdJLTihbBMAnLHWowMVKTX
bM4yIxB/vvL1mSBYjpQKC7o4Llc5dUiPQW5nrdF3zJvSgJsKG6Nt+DCEAV/W1+bTMV4KkJ7VHRCp
Dmida4cQTMxMllZLiUiDhHcsDcL1UCR2T4kwdYkQ+jdnZKkPmbbZmMF/kMx0tT/3KATOf6jEMyTY
o2obxSUxrRzqr/0cvQAxYe+d1O22MbCci5GRXyJhqIY1qiFRbEb7HRyMD9NUGQEPmx18CuJDTDUH
twmSSXNXuIPYKIPfU15EsckpmyEeKybIWILpJoDLasrB7uKBcyDf834kdXpbrRIhk+89DbI6zHlo
1Lg4xadtHc2JfHwtPOZKlf7EFZNKeu14r7zetsgxxw/ZqS+XYcsH+TKE+yYl6yS0Q+/GFe+wAD5Q
bG0sEWA9DGLaGaATWOWC72ZL9QkGACIs2P+PRdY/8ktiEYqyXf9SoyBhOftVcw6EnfPfG/nv4akK
rjboYkBckabPp2cuKguSJrbwwAHsbyI7ZabUJ1G567FL/fjymBScCpomlw/SmfqOvk7DP/ji/VsR
SBiouMOhCddy1AJNoTc+jnCM+lSdDaHxSj2zn3gnP+arxcVLqC5fWjk6mx5WkvQsE1DziE2KpbGz
mT9/osnEGI5wZ+mfICsZIpD1Az8ESVt0G4j7CrSebB6FoWMRVHmAXC/Dyyf2t6M9bT3wzRRffOoI
Os3DgvVSBGueJ0gf/e3GxOgR03oC+4J3NEfh8kVFTIg1r2/UomksgGggDDqfM7J9ftiN0o4SS2kc
mEIlP9fWKJ5au1DfKzcMp3emMkAT27HRkK8pM/Qv8gRm5bMduL/ifSJHXVkrTqe5xIeYjJwwbVZo
+A1ZxqROYVpnJ1gC2chz07xXAdabworEI+JfrIm+KkO4S0XRGu9LjZM8XB5qCn+nUu0inLzzyBDv
WAXCgTdI0oZ2Ef+NgjVABGk8VYfL9TqtvdkS9gCXptn6OLiK4smfrbJn6t7kyefEdpnYggQIzyWm
hdO3x85p2ZTCwxahzl7dFU7/WCofshzxzO1qLZ8E0WC8yE4DMbnQHUuPoA+q3I+njNZAeTRfrVsK
SPKHHugIvZykAuztg5Atd1q46BqSaoWzhOWz7H4QANdy2fS3w9nMAxDXL9+iF0VxJNMMih53ZB+c
AZbN0wWxQKahUah2BO89bBCekvkghI9v1Lwvcxh0shI2Ua7zczL41i589DUbuMEjSTElsoG4lCZe
KrDGru5eCAhQRGh92RtgLXvk2wiEhyHPV0V/Os64vj39X7l2Xer5QLuaozHpDQ+aUnI++RZJipFj
6sKxfyBCZbV7ZB4bpLxPlDTtpGM1peDyJdJR3IkwMj6nOZYZ/WpGTcFND9O6LZusiNeAyPlg99C5
oK6Ld96v+8wCSlLn9HhV8UoIWREyju6uqJy6mCwrxK1m50QnWUeXLIe5r6HAZ7IwploTnWiAjwCP
TVk+GufnqXN4RbUTZaxn6SI8603/w11yPUUEesax8NZdtyj8iS0MxztA4x7Boz3EM3JRWFCVGfTV
d0MoWDD0Lpqlf7lEZdkShVmN4DClEKpVbEEQ4gR7uTuDTT6oTG+gNL/9oTKjNM4G1rF4aZnaLtXA
/KYgX+rjtQLx6hCdVuXVOl9FJC1M+II0rhOltORMjL0l1Nj5uWLeW7k+nOd2EDkrJX8G9TWL727l
rjoR4FQ8X3IBJ2tdQL+II8zdE0A+Q5xU+j77pJNEyz5ho05yowexcCKnGg1yOB+cefGCMVeXuNad
2cs5gVxCgYVAqyCruNTvD+k/A9zwDGvcKEfzMupy1OJHp9Y0Jbop0f5osBT76FOXF70avwhEbBoO
UCvDKpOntpgiTVXSzBnjPUDviaYYzmRjC2TRnyW7wDvvKhBSX/83HGvX1cwTgthcsUOYDg7RzEbI
t1iQOTCnQvh19q4nuxMN+89B3Pwq0Y63+0+eO4ggaPigYhcx8QUjmIpKeVVJhz7WcWEYJYcGoM5H
6zdof75ffRC9Wnk6l4b7Tsu9CVBsgJaFFJhk/QYpALyrIwRHBYYroJ9Mna0BYBez3kLZ4+zE5Ygc
KjX5TLrpeF9OBesC/iI4gk+9dBZ9ag+PupGlavE2z7HK7jQnfiBe9hBuSHy2vTHHF85km/hvTMSi
pt2Dh3ulG8uJ6+qKi66mtL26bH3BddxFUNPpDeYVnz+q3cJDWuI4HNyrWnSrb29D2Y8FYcM8iZ5X
I9j0RO+skaQ6mcCpnsGF8iFAhhRp7jCombXKSQzZjD5G71D4mLLdAeyVi2Ip1hWh+qrqeN0MxQpf
Z3wKfVZhhNJrXe66iKlc6YmDhupKkMOTdcNLuAhThq3VPYPAuAd89sgHTVslTuY9EESsJ67d024B
IN+gu2EWqT4cvumIzIo/q460LIP5atlcuptPpyjgd5mCOYlh3apGdagNrdlbaI8AhzT50lfqdqzx
r++WIYNYk/NCiasvEqYQDix9myrGEtOqIn2GTleSrDkCSANEDl9vrRY+AmCyreQusJuwTMqWway0
Mkx6m8GwVQaneA42hH7VQ6c3FclBFZ9CDDU3nA5sPXdEfmUn2BBVLu2YHGjFtZqxJ9/oXrNYxZ7W
wdhLtz7Z9E/N8V+cL5DEQqd0vCwU3VJipbcMh7KDsCCb+jFqQxXbG6vDMPp36g+zQsDgiLF6Vrdl
lCcFGdTVZOrkiRME6gRZ+DFY6Efw8FCZLrWONAqlp3EBfujj7DY6YvK9NKOirDQVQoQnahc5F/IM
nLMES+V8xJp51r1TcUTQHDxTcWA/xhysdv2anJF3svG7Gljygn2t3dwkd8SbYSbzknZWfF2sE792
dZ6sTscEmdEcrXo3AsOhJsw4DOr4a9vWwTbXHDfAfYRdjU84d0Ww28Q2j98krVDKtMrx6+OvIngf
wtUe0m8Qc1sVe4SyzN6x1v5e1onWtR66xmUlE7j/LrmjKWeeb3NToI20s9wln5ZGEebdMAY6vEbf
xoBrwDpUN/K8QWEdhbtxmaij2kj7DcarJYRvemcLs5SdKg9ZIJt8l+pd2MQCTiHUa+GJZWLWhTst
W9lQq8agj8szpIj/L7pXYKodYoCjKKjBr0M2DXf4qZnUdDYfOJ582KHzMCA2sysnJfKAQxn2MfG/
IS8woeBpfus2Zks940NpldI3HgWgIKcM9U3BXv45jSXhqQkoGUqI20BYTMyS0kj3AGksvyedPtAi
+bdhuiJSJsP/hFnOs9jo1PQZbHv7vtJkdizrMwYDrn5MgRsSUwGJtkBA6IMFvCFqnuoFYOeeT7gY
EUrP4lWgJm9WdZGizyHtTpb0Fvpl0jDhHtm4kiDrJ5U5YWVoFyhLKMyuDpwGe5OZfH/w9CiWHzhX
nhmG2g551ZRUM1sum11DKL1r5nK41HPlq4RkNarkkXAYwl2WERipUZ5m9btGI8PPhYr4wDmF6Ioc
XzcqocQeCcWiJRjnNK6bxlt5NKbUHL0/Y/W/V9W/AYLRkFA4naLVICsoLyvHWUTHNy2FQxJq4rCe
Cn9IHrfpJsZDDKRt9nwDVYGIBNwxXy6LduY8vjPGg7ZPPhOGe2CEz1YdrydBAsJldhdUlGzrJYJE
gizF6ZGwi5nG3fOuvm8ZRMkEmJw40szcqfN/SrWdQi3OyP8pYBIQBMsg0Nkwgq5YaWM/017g22qT
DdUpcJl3fg/v7I/l66iiZT+BxKXA/gkpj4rgLBwt2yzyn7TZv0qF8ficCP28KH9ykMupyu6D+6N+
gM3nA4H97ck962RHCMXCuMQ2Lyz/z9AbKNRhP4nXbSlUJl2cPcejfbwqJAWfaWrS9Uj5kjMJbt7r
tSs5n4KJld1ItYPKdql2JBln0ZuN6HfkUVaWMp9AliRqIfbgCWSgeaz+A/qcAOUBKmm+K+ns1LCd
CoHx4px2suE5o670EWQ7BohTbvxKNsbWLJdEymhW/5V2EyO7zO/FzkMlIuptfO8hKh0AXg8i6x3h
/+6shZJo5CPIyNCeLIc7bmdbCrcvDWLseC0s397szOYhqfEhD+EXcetd7wUVZ9Pq0SPFbesmDndK
A9moJgWPtK4stJuTu9Isk3rxPeruJPDMt13kMk3ooA3DzxtxUtn5oBKK3szx9uc90835TRJGspVw
HVK/zSfcuC7OibGdcCkhHLoTBJtVy6Oj/MKPLB4MY+yS7X84cbugIRlt5bZyn08g80vVH6O2n0Ct
Xo5YVxmp7HCoKz9sGdWmEBqFOIQTJ7OW9KvpcdflUtifMzOiVyhzEZvlW8ZsBSLyf9ejgsIjePzy
F7yfwvjlFdcaSG6DSn54aYhAhVkmIB+TJQAJPJUwqlf6vHi4GzTe/XDgcnjV/tW85IcGDmXJ5fSw
Js1dFF0B3pLGbo6kwwXk3ukJEcgBxSGYSbnkJsG4sqSUQpQIgeeEWooD0G7KjFDd5SFoNMuciUcr
2PQxEXLSgFrinG3w+4W5urrTlw9lE9aw3RS4SJXZ/jRTknHIfd8UpqxqoWOHBrgAjWWlVF3OHnqo
kgrwPDkUyItk3M574UoJFwFzsQI2KFOZE0yVWalUtMht20O3+65XLtqMITSjJ3GlcNKYqmwhu1cV
f+OHV956n1DAlVUxTiKz3QfeWpXtv/RTNwJrzSdhv0zgmiBGfVL+3ajApL/T5vIudGArAMga+Tf6
scXJ1PzdFclSl3XFlrIKkmWq3Dwv4S7ct/tKVAfNHDrhAFeO+mJZmdltC/eyVZKdQLv61ONVbmx4
dJeI51ez2YKcyRMhYa/bYggQhu2ZhujZjPPFIs5XQCfDrmm/WlhLYOagGA1yGgOd3ZPYK0BCs8+H
wIKW6X+QXDz6+L+t+Hreaqgq6MwhsfdkoSWOYCTi1/BqHjSWMNiaqgusiMHVlUhoLj7XNhwks79j
XuaDs1sVnH7+719rdHT8nqws1rxYeRBbeHr6c+u5BoXFj6aDikZYxMKW6C4a05gAx8Iwtps/qHQf
fZtl/7P5T4fo0L8VYj7MGCZat/+h+/kYSjnfm/6A/mDxvuWzwSal1QP0pS4L9DCiEO6KH0C0WXDh
fNAhBUfYYLUZZIjPgnDARNRu73+DvWRrGyrziOBYyZhrAkbpnMKuCvSYIdbZijWQ34Jq/zV1WXmN
JA45Ns1XxRhbzoyQMxw3nGLlYbyGfmrcmZYE5lwDnSoZKSJL/1oOldHjs5jE//A7sqb+3+Xia5Qc
UP17K4zQ9Pi7MjLrwkZSbGZuCtK5wwNDAwYEyq6B/4lyevMcq0/3JbVqJgXHqfT4FVUGR605LA83
sVLVTpzql0GgaNQem77nKYS3mNwp8c05d6Or1v6GFZ+NHLLuE4ujhlwfmUM4ZrIb7C6Ld0njW/5H
xM9S09FUzJn9j78GRONv6c1CrC3v55FVNn65NyThG00oWNWMHepbf6de/LQHD6O7/ZxdeZKYT6ih
gvdOn7OtatIiDH4ctQ4NcP0Ms2RMa1GIhl1nKidX0U6uEc+ajXbkK77Iz22AOOsQATuTFG/oIrOQ
QsNBwe0MBHKtDdKjGqPOtqqkfmKnFlyH6MvF/LfHDz96dWyBRuKnZ2mbU4+qw5qmDrbxYPyTXdDO
qiVF2z47zZQ1GYp3Pn5Jlm6vNdogL5iMTq/6a3lK70r7I13jVmBr44K2I5LPy8fU+FSGjqcHNSSo
1c0hsx1xuTDX8Wid7RqZ8Qz7ThjsMdmsQA9GjMENw7JY1zJettecek8MA+cjUGpcJ34wBh6d3YeP
iuIGWAZfw/TZ9fmvumNY/xxet8OyFpkU5+xCfOLLeiesoqz7kPCOBQN6MQShlVkCED05WfmFx/9D
EeWeO0MYvJ6OLtenCVrxfJiA8BJ7rxVpz+5aPwv8stMAiTSwBLBn7cuJNa0Z8wTOI9f1dseLNfe2
Q0d8MxhN63uZDamQp8tmVEtYt6ccV3S31ZNozsJKULHqXlBqJncIh9YX3D9YUdssTY50b2SpyxOg
weZE/iTfOeC04qUccUg36j1BwIlNHuzT70FPXLx8i3C8vKnKbr81ebNI/GoKN1ljgWEXtrmrmszW
wbFb+SCMh92Gq4m98TrQ2OU0qHYo8zq6Fbhfc3JPY4/2pttnBfvmbzMrs0BcIW0jdAmjN/nsh7Ne
uZ6Iqp+jD4vJWoEdxM8gba+f1b+yrdB5KL3qI18DEAvHDdC26ydePlVYZjv3z6hOnOsufcqcRLiJ
FrWCagoMlb9tLMu6nf1mY5bX3I5aXkhMppTaQaM07f/EA2XcSE9sDBQk1XkU1o4rmjq+ld/G7whP
d0I889+n6/4Uutol3rUzadY9H7mlEwWomLRCHI29uqk7LnvqpSO75/gxA6JvvFwIl0tBSz/d7zAz
dpZ5zFFuG4C4cDhfOqt6P5Cdhg4arqHScbt1TqxU8jXbgej6Ojqc9U48lgVpqnMM+Ab3DJ4dYZb7
Wtzn/Rmb5pWXYryZnlBJsiLqiuILK6p2G3VzXL48VkG3iqlZsn9T+HQwMBJOiSe9xZ63veFAK17T
rarv14KZ/2VnvC8VvjBymb7+GudELUjpitlxNY2MTO61PFGgSNdwVcudbJYiBAJ+okKyO/e6/krr
P1jK6iq0Y+PLaZZ2X6Jh8jCRwlF8QeZZJcCD1qhFEa/MOsF3tc+ptvsnIaAIj6ZHrKmor42zy1fi
FDGOmvFO3wz1wNzCef5HT+mLpXLEwf1RO8ZnIqkXiaWNpNhvxjKxlG1TY33Ef/KDR5PV+GLDKMZ4
ih2BmnSeUnxQqx3T+nJ/aZ6OEaomSXy2mHyIsOqywJ/9GxJJ0w3MCqiiMrTUMxJ55lp36JAbuqby
98Poyx8oyXEVTeee/1DBut+tvPS1KNMBCjAIOCBxwSPUgovRZ7tBTTooT7jb8kAdBB+rrRYmmCro
WtfRczIfonB+SPfXE02ShPVfywlhYPH322vzvxUKWf52b/dfrTfoker+2T23tvLjPT6/04VBPkN0
DrXYmZpXV914N75E9ROHQGdpK2UDEN2U+KM+A5VQiZVulFWbKOvjF4tsoE14kMeYnd0otQY2aWB4
T9/oYfP1ShGAk3d13iDsTr6zVDlK4MQZRfv0m0ixGW0TMfpgFSbRSaFi2JJTdLzRtA8toNjQu1Wf
ocQErQ0Bis3GXvzoIzt1NIt//kyS9Kb08wGpS60onYun7E8oC8fTg9aXOFuQqt/vFUEPLpx6no57
RuPz35pGnSOJD0CzoflSwGYNq446JefSWBLsWCmI7kqM62+W3i0Jdtb8B2XSFvSA47n6061TwnOO
itDEbCQo5pBnWsG1qVABkU5dotqVCus4P6mVEPCkRg98k21PEn1Yx7Z4ugoQswALGqul3agAE/C/
1xByVfpOULU4B/5kMQVsbCLSYNmWPN0Slh3m142jPjO/cjMnDquORUMWO4nwMcM2VCbelf2mWO9g
4F2QypAZcXx6GH091uOJY+R4dv0q6kiD2rqJZX8SVh979aTuAi3VjJTlmZxvFZpwsFC9g6gUHOOu
NGJue/uoELjAUNwUwQsfdiC+5sMPz+/umR8nJwmtM7om3PyYBPX9WA9YIS8kWVriZnoYgEzlw12f
3mv/9vF/jdTs6WzGeuRvRnyYyQt32kQl4vmTupHEn2wY9M3h0W8ChxRPofHOVjEpX4GGkrCQM1xS
F1rcd9PXo5IjfY6MjSzWoDMpc27nlgsSJXw3wyZ5DplntbeN5wVjeQkGm2zNBgq9Zx07yPRtRjQN
TdO0Db+JWxRscv6u01cThI612/qCMKyxNRXavpuDt36vlIZanjZTUCF8wKK7rdLkVloUYZ+qnGSM
8l9Xtfpp8wim6/8WjScBZ2k3Ul65Vr/7exxmNF6IbsFHjuZsEkSrPwt719mvfeI1vW+dZ75JOAYC
0FScdLOP7g4O1J9y5qtrwn4okg+5UzIwVTW3/8jf/ze0YQ83GpdJEIZ5VvFay/7tfUlbfzHjqpbg
fvrcE2/fQ7w0UoYK0SlZFFnreMBPPvDbRhy0qeFZutGbflJY2rwTcaaGpil+LKdvftQBUsgygZLd
VpVdYNovJjl3sPpbBVz2ieOuI7WSucrTBHsiquj3oM6zDFCQtimKyHQPiN7Y/UBc6MkwmAH5qa4M
lrp4nsegy1mXdR6txa+TMhsskP8l3b1BKVdTXGifM3OClHI7b4FR4OR7BWh3G+ClhxlpTFCnTvSb
5VcGFmfYZOWJsqbqBWbz66+466aHjHu4/Dz3tvOEq3U3VHvJsmT0tLTJwYKdVxcmkXFwOfsuPcV/
DM8tXpvB4svnkN3/EalcHaQaKEH4S2DlshGywzKV1jWNwjyTdwe1yVrkmduUq8ew2agRLK6VW3mM
75zyzRefJCc/oJhbAo+XXdGlJOUsgAVX4cwKUGF5Qahkk/qrtITt9a6E+/14Z3YRs/Mw0M24JEZd
SZSeRjW+Bjf/G6U/axj7z4JnkCOYzlZnZhBF6sD6NWMC+K8MUhbZumikiLWIEAy0mpwVjnuA1U86
nhM/GHaXkQcV3u9R5Ufyp8MU+Zy3pVyatw35r7Mk7crKU685IsNIV2eNxK6XjgD++4wNE+/J85Tg
7Hk1hkXyjjZvEwr72+J/Jx5idKPbaLCZww5n0DU/+zIQ8HNin/mPS/gUSHgwtIApDl6inYDWmCPo
7Hse+usYz3OIbcQ29WGlwAksdbhwXBAvul6dnqozi7bfzHdZsYZMUpqR2XZv4qxvtaXBuKk94wPu
lqjvY1iWNEhlric9MHG6GYQf9D62l/Kg4aeF69tIN8JAT1eKqm222kLofjekUpteJi1hUu/HlwD8
E4tYUE0cMhmQYVRz7hvxULSFAGtfy2YLEqx4bis5RYmzs6WRj4y/deo/PBLGbiD5ScU6ZgTtebHZ
YWzr1BH4fgv+oryXPd+88wC/IOh2HmWikmdCfhkpztDLR0TK9ehr1x7kqlL2ts8zzdQvEwY9dAQp
t0FzIGouyvA0Z3b3W8zFOoGlB2zpsKUUYCo8GWqvKoLBO8qvReLBlgXAPQSFSHGunc3hU34E8FYO
/dk9GG7YNEPwI4Hky2YyWbsVL53QDLtWFqLVhQC4lwArB+XY/zJ2cR95IOT3yj5CoGEt16aUQKLy
PNChxpcA0NrZgRdWXCbEcOTLQDFXQwrR97P0lSo76RWpo9Fy2yQ7PyrLbhihL/7iXGrZ9sKNY4Eg
mdgtym9YRLfFnP84EFD1N5j8R3sC8Xe4I/SPvaYDV4ruurrSIRHJlYmF1hT/dthrDaTpGMuiYKx/
aQQHxkx6NdENm1Sx/QjIZOFVNUCSV/YXI2rwNAP5Ug8t8ptRrribEnR5Ad96RYXf+ledaSrEzIin
ziMGz0S3D+l5KB4Wu4RhcY+yfHzYDDC3ODCgct3bDy5Rn7NPRwtvf5c7uux72zHvuRUSsLgh5rlE
CWbovfwnp7BfSbpSGYm3xkH5ZFpNRJJ6lAJFUAxjyxwJXm3hRuurdTR338Jj/UifICyO7eKkhRWQ
RR6vNjZr8b+ykasD1cSSWBJL3RoHctYBw6Lxz+mpMDXM585YZtydyVpDvi6Fd3EsYYO+shGQ6ut+
WrWOzM5spFlzFGJ1gNjx7EcDQSrNeV0rPU3ExsYJ93+/sbEIGz82lQqM0234yEtbcKCQ6gnJ86z9
W8xcOMq57XmHu8VUYgbRmrSY4X6AxsdA5q1MFYlQtyEribVeidDFakGykPreCBRaawTbjpuQmaI3
8Dix/TTKS0L+FTrXPeiWg/z2D/s4IliJ6DCZn+ds3VMFZqoE9FULReVU6Nsk/ltLVf+xkV4kqY4r
LJ8eBAENu1CGHlG26T5p36oMVpcnQnGvNqk03AWUbemfFh81yYWeXj9bERftCiCqbulxZX1zefo9
n7jWHgOkmgwYeK/F56jozW2cGVMv1qeZkLYXpNtYmrUa/TAANK+YBnPmAqEzywSbfaftaMSmrFbA
8IB4UOHZ+lcOvvycnV5xLXSy5HpNCBq1stGZc9FChUdzGJ+N6SJeo1Su/FlvI4TotIy1/FzrnL87
trGMTZvOste2lFVAAgskO4rYVTmDQfFxBnWhF0YT26lv5/UBftac0CVNjtkEueHwX00tFKqKgzUb
XLsLvDU9uDiSG/rcc3yiBWho/AcgtQM5n+bO8CK1UXnlJBicZlXZHHZtb55NpodE2OL5n06f3fWi
A3z7LBBf6xpdjUPCJcUD5RWy2md/cAeHBZgC895x8E5US5dZ+VkiTLj3ppEIfAiXhiMX0E6tX3hd
/dks2kyq6n3aOYOqe0A2hzjY7gHuXQO0B0Xy5nM/Dhk6Fd+CLB2yutOKkSseSB3HGFBM/+i/5J8F
zinhfm6lgNOZZRB7il/GZn54GL15G5Dx+0/gIHCaSIw/Z06JAAjNLnMLU/8fIFsW5DYve5w3gf+Y
6AJTyOzlcZ51JVDswRh2yEtmb9qMImFZsfgP6C205MssQApHv4LJ0lTb1iADT3h/bOFiIKUngD5Z
MUVBjb7EO7zIykBwWyx+vj9bKHRkdzX/+vo90NvZLkresElonpuyXc0gvHFnJORsHiTDjcXc/XDI
/ml4DzM4ePT2X1QqZ8NJ3s2B9vVFLCmDNyLbu/S3mhD2wNJrHxHplrBERYUvz1kd9YBUTkPOuvVw
QzS568GuvKGog2rFgT1JNrIX/quY7++P3QgNegW2BNdkMYOtUJ67HU5hxZD+dSWCTYO95u/Zu7oU
uf6Qg/SoPTOhaqYpkLLJ4GXe2hyANrF+Txw/rUdYXuC4rEjJ+5UfdX652b31w1Ytx1NvKNRq4wYI
OJvcvAb3C5+qKgIPF3sx0JHEhYbxDAd/tHPWuhLtySmk+1OGH2dZ5utuIRto5ZecGISoHLxZCX9f
4XbqyQdPj7yFOa6HC4xlCbU6YkDjKzEV47sFgTOxvPmBezlhD7dT5DZBfSQQu6PDPuAUON+WqsdA
+L/yo7wEbRaJghFMzoOItb7bgNvjTtjFLABlWUwwI08uRjwsA8YmiqiJaFNlGqlYqFZL5TSZbXjU
XTc5dXQwGgCTK7AZccw7FRd/zpdIy5nGEcPUh01Ol8P4ln+HLGuZKeqYFyMv8aEt22nfS7osXVYp
mlUnYC6Wlog1krErdh1okIuBG/wLeqwgjHbpPNC75p0y86p8KB5hc1nnFRuVK2hElo4/3h+N0i+k
qtQflvZeLZpab5JK6YIKbQoAylJviu4tcst3Q7odEp1qHF1ePhzRkqhydyEnokVkYnSMryf07YQN
0BQR0nPKGPjcoxHXkSEp5vzzV3jNc4B6qP2eOO0b2N5/juCEjsa1s58ZOaoK6U2dj9Vzp0NH8aYv
nse0aJ8sGFT8A6z5wiuSDPI2s34i2ocS5bJS5baX1UyggpFdgrrS7K0N0OJzLhwktRxD81mZGf0V
NZofCC0mByraZbV6BNKTo6NqhEFiXD+8GO6uiucsJ/18/kKujxwgOtmCkYMsyzkmmrQA3Qiwa+1M
Nx8cQY/NZD6OO122GTPTpux+hdqOJgKV9HXFgUblCdepSnwc/wtNzD4qVxYBpqYSn9lVluZphgAk
NfFYFGKYDO/fKaoU68OY8+BL/DGKOF3304V54kpfD+5qWJRk4iDtrEj9ElMHgvkudu67l0+NmNRV
TW6yheoXaSG6k/4CBqLzfs+wQrl5nuI0SGsGZjpO2GmrgylQ3/j5Pmc1AgmkjIrI3NpSQo6h4ef/
qEw4627lP39zlkrPCGkHmRx4NKa9npLxysmEJAOmmArwRoTjQ7W53k81MRtdHYtDaWv+bUN7FqWC
zeUzYL9KciEHAM2jFqIIJrNjitSEhk90d99K2WNKcFYn0++BDa/semPVMm2sewfXlsA9uQ2DOtsk
/73CJ9A7GBhyrb5q36KIKmVLOa5t3LgjXIOMSxZy8X41t82h7nwuKJO57JKhnVj+jN9NlwG6fJAf
x6M18JdQ2lGvLILy154QXciR72O6K6jjlQyOee5sWdipA41D3wDdUDtn9FpOYIKtLkjudv4KIjVW
eOrQfqEEpMEaPKfNdYIUzz4Q0HRbphaEg6K+tECyhai04fFt54FBrl8BCNwLYgP0vivuMo2XUWye
o7LVNehtjNy4tFhlDEqLacmANQiflwFddfb/agrzoan2XMb3NxBR0QmgazGu1xm+7NszHv0h1aVI
efE96NZRcV1N+vhOjMQqVzx6gRpqTPB+6YIpEeeD2rNMwvueqnCz0UwA9AljBI4pTxb0Qc5yd8Wb
Lgfvit0PJx0wGmD2gmuMmJDxfR4RDXWRo5BFQ2p26nkQvopTcI/YzHdNWjWhIci+46h5fl1aOz/Q
tTwtWdKNK6qdjpNRvTWQXaYr/K6dgZGFQ8u0Ha5mvcgE8ZOwoa6V3Dsn8KjJaS/HgW+/57jVCLR4
eGd9ADThlv6JTgdXAKpRglSp3JBuzZXtVhXPiv9cjPZL8/sS83JTbMEfg4dCi++dxLNA5wzIHDBX
CaI95PUOixhCmoFHFfZIFRoEIcBH/O2xLbSFXpoXIeoRtCgZ78+f349VsGWvQnUO5Y/orKwBY4Ry
Ab9mAERA29WK9KZ8N92WIpf12NkEBko2sef7MbPIqfWcjbtvoNWqGtn2XUfGimkIAfMDA49VkBUP
x0KlcqmGBkjCKnzULKLlQeYG5I6NgsZUZOSVXB+TgvCJYV7IkkcY6nB03W+o3KG5B+x00trhBDDq
DCvJoJ/KqyNgtH3w9S0FWLWctNWbDTfDMeHcl9k3FR5119Pbjxu/w/m4NLD7pnA69MgD1tt71YPt
ZdORizbE5zvVPK8yVTbgXDfBJ26cMHQFOm6LqL87ADBgH7S4bN+oCWcSsPlTOEzObZUDjJDx7Xzg
BaT6i6pd9cS/VZKisAyKC5Z8Vgi6kjoen9JEYXmOOS7DH6d9wrDZABCPQtAmPBRdoVT3jt8BgAgw
oT/SqTFlMI11yn4mbPDX1Pt18bGBo9jZN7VNwI8slQpDDoJibEcTCcUvIjsK7J14hnvJaLYRVkAa
7eQT8DpLhS2u3TY8Il/GYFqY0I4zg7dPjKPF9fnQFAQuZD9WI6R6q9uBzoc+4jvRM5BmKWLB7vBg
7c6kgMM8ZztSb2my50qlj+3PuMMYCiQ+3ff6iGit70YRWghUoUHJMM/gozw9U5dLBOPNcSBC0Evq
zAPD5yVWe2eUjty4vDhJ5EMzOP50IA6A9B8bFQH6sWNH4yApcubBHr7aVkBLIywSkHi2HIAGKmgP
oWuiYb3xPVTpFX2Yn2c4bJco+k7liiEFfsq5GHUDQLFix2+2aLMIZBrZLwDGjAdUzsM/ZBFyATPo
pgYS9FYvRvWu1FbkW80AXckuxJnVPcD8mGqUz6fhp+ZgIAEi5jvn4XCOfk05jXG9/g0JwDf8uYH0
Gke3B/Oyk1Qe8b8hfA/KPLIUGxQlYBr1hHYZIGeHeCp6gi79zqWd1DLMvoY4ycLH9RUG74H/v0Ex
cMreKcfeRW5wJqtHKv/r5WhcfuhW+OognEgPzw5n6nl6oQ+PkRJ8QEdByb2plOiSJuydcQkLQuo6
aVKaBZlnu6Of583zkezPOtawrQ1hF8lT4jnXCRZMm+KxHhx9DgFtxjvV6aoQYrVmHb5cg86SUxtT
mUYk5VYN2gb7OOfd5+e/oE6Erz4E+4iY3TiF9nJP480J/ucBXSgBklPsaD4w9WYH5N238lFdY7b4
YIvN0IurH8iokpPozgxyXmEVtHLx2dFKdcTsKQ3gJBMQPrHfEZuZsqLgNyDkt2bhP/Ji/9MBgI4w
AeemgriASwDTdf1A0UCSaTlVYzbcDeEEifOzLzwDDTTVwj+6OGoBAT3ySx8dx2HxJ+BknT2VJYSp
BDQPOt24vadHYUYWfYb92RpRMnDK3LdsP8zYkr5szIpu964xDtKA6xZVUWbgdsxcBG7P8PmvMlzR
NNGk96X7KDNzANCOtYwB5PWYwjJs/NejWE7z6SIrdy69FMMY2jUOanTsTBMgaP6PKW28/qqO5Cqv
HYzyRQHxEIpcV+2VsgexQyWjWjxf0Xzhczf/+hxIU3YO65Gwd1f8PTHFE12Yfozf2UygtTQW7HBg
E+27rXB0c1lCDwwHtf0WaDGiizcu9Rw75eq012mOMx5ChqV4pGvt5v7Akpv9K8AIP4u5LrKJs0/C
BMqHJ/L5gMKVcRSyafoF//dVe00UNRO/jpMazg2zh5LJSXqh/0toMbabQHloajc1Rt9zYIsXEhFb
Tz2FElYYUXoI+OIoDuErb4RMZs+Q8oPywKXUqjDPfPuvorAcNfjYEXd+VuSiPMO8fPBa3nYDIEdW
Bkb6jZBlqVNz0BQuEBPlqepA6TCjaJy1aLjMirjwg/OlIelTaRXq5fAeHaCXtFLZMDW7nayZxb9m
SpOa9vVOJL8G1O/lcDv/GKsPNax1Kapy3FR+TiQvSb5UwRC1uEJ66aC386yi8aihqzGOG1O80WS5
wZkKl2cPSJb4TlbY1YeigAK+ZD/3jO2xhHp0I7FTU/3ekNXwOp1lBnsxg1nlPfppxdfp0eTi3w7F
u/TamUHMvSra2HibMAmyqTtszlFYUtwRVJo7K29y7TFcEw2spfXZmZnUBYkR+eT55TVsP7vasU9p
spDx23zSgISKZOpl7ioECcHwN205cdWQHycnlaTcPEQQD8eZDaRJ27dpbFUaeUpxLk897+02NslC
EspHskCNy3yC4ocNVtagKS9Mwj5ZbwwUZ63318R1IHwb1i0ZZ0GRBz5s2AjJGSSJi4nQKU0vmic1
AtTz0p04Xa7n/9hEMRqNugrx6g0FKz+v9G036TSpdNWZ0p9i9dqJtqxZ0s50Njp90jIXRii8kyAX
MG426CV+KfR9j4yBjNDNJdKnFh3LG4iGUHo7J5HUpqSHLPqGkLLsXsI8rlrijubIT77L3PMVpH1L
mBGMEjcNNK9PvQR1GfthW7Rr5YheZ2p3pRkBau+/da8nCnt+Bxlq7Ky6AzlUdM234mzFLhb0Blz0
Kh6UNt6q39z2LdlAG7oZ4rU2FxgFrjixVAx1o3kO272BG2UZBfpf7Ysts1VGCAu7i1cJYENwaqDY
8FCWAUzJHYWWTFbEP/Hpa6ZyKeTdGgWhN5OYqeFJ3fPMw5ld6BkXHqOqdtFneFVpdBqPEZ4mmhio
gDDoC95wd5rjT6SElHwAFTU//AZeResXIoB8tj0Bp3PY3Few/SeozGjvrcAWlZ6Qf7PORMh4gEOs
SPiU6InW6WXLDAudm5VoTL4QXIB37NNhKXcLNgG0kSfrRuEenEm74Odg7sFJ1KsVdoABLpVkjmoC
uh1bblZMMlGzUjnz/53Wx+z+E48vcnBYU6H1hyMFIcZ9PqcK5JYQYqpitdGQMJRAgYKQHi59Q2jT
UaEZvW+n9e1R8skb1Jg+fRIJmnWpT8GkRDIcnGoD4Qh1H36sWybm36kOsqxOkW11A5mkMXrbAj46
VGoWb9FZFvbPKlOPd38wm8Pnw7tqdXS4NDzhZrUpufPr/LY08wwQR8dmE91CujrPBH5EUze7tlLO
Ny83oAmmYPs/JxoI80BpSi2CNRF8t2P8nEZcPpwbTGbtbn/B9pc1r3dL2WcxVAC006lWpxRYzG8E
q3OiIIJbJ2uUbNwxeyxkLuOO+gWvQww4D80ADSw8CwK0QNDuJWciiwjfL17VfOcxck//VBOo9CnG
lVvOcU4PUMSSyVVss9k3d/AtUOZXbX25h2kxcyXPbH8G9h9Z1IqWwYN27NtH0hH8MHgsgPTEmZ4w
YoUIRBKUwQXpIhaSmIyMwpofrQywQNaqAOO2OaRf80rX6JI/WDioY0gUCxo0wno7tfZpKuKqgUru
M8nSic40q6LVfRjk2BoGOd/nfPZlauWumnCzzjrFKyTQDCwf1wXGJKkXLWA7u6txmkJ8LNafACqc
7+hDss6/ySqsZdtCnrwp2U30c5yUJACevmrqn8k9cK/VkxpQZsykJruzaHiv+aGZt5lrhhr+uce+
fhtpRveVdv5L7TB2gMr5hymw2otHh4s3+rAi9Qz1ed7Le88JcZA/iiDpXwOsU+RX2lM0neRTL+bd
OiGnr5bNqoVlWIFbAzZL6yLHFVafl3ceL5I90hK8vUPWOJDsz4cwdc6LbuO8na1h8a2rEirJp4zR
41nt3+dZH7lN+dZqr3icysPXzpw8Q58YMjXAiDk3mmdaY6Jo90q6O0Sy1BjNxYjViwpu7suQzOt9
zhv/4aNaabyEYIHT06kdLdOS7a2yswohd32dOXckEca4SdSLMUirU8WLIqvXdMUA5y+i0kpKXuzy
C4WQEg8AUrQ5wqQE0dDo/q9ihPMEVItCP61ZYTXjRiTM1j/ZtpfySh/W9riND6XeMwtdcN/J5ram
nlNGtNeKcOnB6fGB59eRS+kOkT44WKNquZWwe0Veri31EcnYcwEK78lMF9B0uPp2ETKBRG312zQZ
WRkKQlq/NF71lsUruV6Xj4e+CNyDLRKSdA6PVREFMMVtlqmIlqXYPafRRDozErh9cUNJ2+2OqwZG
hEFoMsg3cULteweshqAemXDzAKW0xF2/eI7b9fEmRITgd0E2pj4m1CwJPuAh1K9SivufaO+2c+Xd
tWYxUYnQg7zsStcC5pEHMgfGkvLQf6cIEis12s7whiu3HWdjbDCuL6HYXO2ZGAGkl/hxpZ9Ge7bI
tI/TwhyowfTE2u6PxL+6QBE70EyrHZwmusIhJ9TOPGNKEXJummPbiiARE5ldi9MO4Lhsn5WlaRQf
K/kZw6NFF6JkLNtiGWSZKMCBnykPgZeXYUw+lPX0Fq/bls60GiAT3AgSnM/bByjIET2GrIa5hP7p
T7AspIj3JeKWhq1BV0srzWZJPgFVnq5fOUZ+vURZw6uGTAvwdH2FJZh2mUf4W/zEICFgR9fGEPRk
A2S7L2+BC81r7eWFGpsMYxuXmZnUC0NCaHGa/5lGG/PROiRjkst2jNf7emXJXR8lW2IUACVSAqHr
HwjuzOrZ16rabaKOCgUgp8TWtR24TEN2vlJGsl0m54vJvkDuOGBnQdOKf/SJCI+16L4wUFK4U+Tn
8kadzQm5pxoqvflHEteiufrRL7gX/xJAPLUx9VuQB32S5W/EN/W3yhdnli8rvmQwxztRjHDOTws+
KfdBK7RofWeIoenc2Gp40bj4IV93/R5IJDCV10OmXW6bGQoSgIp+rCvfML3DPK1pgV2R/xIb2r4W
MpHi+LS1vjuFrgS1BhTDveX+zFr0gQE1bXxzO/N4uKE3NXz5SJKi6SVhJqw0Lr2mia0z7N+E7CKt
AerD4QR+HZoLyds5294xHgpJJeXCmitIM3cV0sfYrdbml32Zkhy7luV4NsaDmL9qVumf3R51v3RQ
y91wADbwCULXEDurRzGXmn+FDtpCb+p8TQcrMm782R+SGSiyNkAjohRvzuypddoz1Ij3+oaP56fe
QrWgD9A7RCd6JO0dOlnJMbkU0iT1sUJSVltl0sZxbtIsOauY+EhoYUd/dEvMJffwttswODFmdzM7
kGk3YfMkUjjYg18p1/5wtIRYKf0kdRv58gC0kLd4Lkgoyv8zUIPbK7YSpTq0Sfat1tIl3/VPQION
L38oA0/GSv8A6DlzyhAmCC5+fYdbT4hKcrWzAqV4rMTS0t6uw3N0NTvlBH0JPsM9UAo9G3TEHqpE
PpEYRcqyUK0CEu+NmcXfVSsxv6HOck59ZJGD2clKFv3AMBcpQsDtzl54VYXwvKfG+ymC5zUUNHp6
uNhGlRekDmbgCSaXf/fEFsOrDHdW73QN3xMpK88trqw3OAqO/KdJ4/JnJuvfnLfGatIPqahrKc7A
visbHoZL8nJYuqK6KLzJ+s6XTYlv2cZeQjqzEN7pjZyC/2jHa2Ul1/TgwegFYKiyL6oFT5g5PTfS
8ccXzNBJLuK7OwVCof5eaO3N+mkgrpoeyMKmmCqoHgTd4IWSF1pudY1tgXVIStyOMgT2oZife0fA
bBtRzBfGpVAQ/CwJs6zo+7/LTgjzd2pJDEE/FJCNpUBs704s8aJURI0shU+W5WTWYtCtzw1A6QJL
ZUtIdPxejlpuEay5uMjIjbxFtS898gIfTbgNIcqgYQcF0OFEO0rRqoGAsLKEvB2ySnqxQvtFtYC5
ROInrh3RA9SjtRaF0TxvIspwbZcYjZUbYUBui25vPx6SdNFP3qIP1yDwf9AUxQQLF2Gt1mkPEYP0
mOAyb+8gp+baR7Uc0VXDIenZf+ra6dVZSXzHvYBGOs3zYCGweakQ8PdRsja5DBZysDpDFIuuNZ5l
sUGJoBFzlX/WmpBWheDdyXjM/cvf+W51rtRriBHKXu8Duua6p9RopckYbtRRBJn9SjCikZcQQg0R
J4tsj7yz8+FV4BZg7JDyZZQao92QYvSnwpYODcQP+MAZLFa32tnC1ITqED5A5KTy8jMLoPAL5/Z7
B4g/PCQMhm212xHbQmSdSpKN9LuUvVVXeZoI4Y/A3ySLqtOJlTzH8Zf8DBAoUGJ8k0jPAV4XGFlo
HFeXX1eB6qBtkOFiNthfxuBG+mE516U6dczQIY6nn41c1p2bWuM2HLktKvxskLttDLHlWk4fdKOg
Et0vYmVlvyGOldKYxyeGXGoJg9MDn5EPQtyKNXSYYLDpeii3yU8nfJeIGYrfBkEHEAYWjiJwc0nb
ZEd5w9fWvQgyCPZ6A7M84i8/aUTuIi2WGmXG2nlZ4dnqZoPOzdv6ISnCknMqNLc/eM1nrfFKpT8A
i/MDQLNxU5K97PiRUo3yoSYJO1SY4dOSmICqP5lTEfU5R3YvM+cX6+PsmmaikSU8YmpfcanG2NLw
WYTlJhRsvISXJF2YNkyI0bBAIeAHfh+OqD4UyNEGr1Iu09fe33DTugCNAm73VX3783S48EUi1K4G
DlG2ny6vPHgBa7wUBfcKyksekkimARCEsudhkGnhGs1cSgVCAnKGjVm+cw+dvRmr1tO1/kkhm1Oe
PD2J5a78wlN4ZiLuRE0Ax1jd5TO8VTm5nCjytE3wfUcjHqmt5gSajrhZ385Cep/Af81BH4bdH5Hh
w7/KjxfgmXOIeUQPvMYqXBh527PEJE//c51V1RtM0M+DEsaQJtSs5D0Ibmotxe6TntebAIqzFP0b
qxR205t1R06FKSH3+gh3Z9QXToxyCrOWvo/SFm8I+ZBKZRYvGGJ8kBIiH8989gk0R5MIJk9qNpAS
FuYrHyAyE6v9YkqPdBIsSdkAK1O1yKLQiIEs0qve8wPlPJ/xMqI7N2PSyJkQWFL8Z9PB3gX8P5/5
Hxhvp5CqYQlcTb4QPT+46LpqfDZyeyQAmtTB9Ed6VMbKEYPpsmwPDfpwaTdnr5vi61U/o3SqAk+N
uBV3YFX4h3KJ9Qa2LsaRsJyk8vVeXfGEUhL0W2fWUBoEB4KGQIxda1vuJoTyEZqsqwulq6554ba9
1XletcbwynNgeD9dqvUBXhZWDAFmv3QSBe2vN+vUodXDrMGQFOJaDQQoBdk68f172n2A3QE3XDPe
ginzfXXi+k0JjZq9Dq6Sst1kD3Wxoo4D+9s160fU9Kho4Ee+2JVXO4G5EhRRpTInX8DyDN+jpnlU
GFwl+hIBds5U39vBv/l3GdYtrsSzqYztkL7DZqE0Nxi/LYInSAqfSEbYPPOeXD3h89wRu/GO38gM
FuK11jbfIpUFgnhIBBJAgAAtpb9n07GnJK/cN+rw+MO6J9AueCLjaAwzl/pMr4INtu1WvsRFQZDW
6FJJsLt00PheaUk+bKdbxWRRPJPwD0M23CI8awWJ6CyeNj9+dpnI1FgVMK2CjA40JPHn2LkA+JKR
XKV7eAlSCrNT8SxwzmW+KGKb+8D8spm12lo1YTxLHReWCUu0vBVCUiTq6eiaeF3pNxDOQRkEWLkw
bBQt/wIJNKrjDt7t9CSQ20VfFbLa/gJ+JfsVGuId0/BM/P3iRLiH5VJBmojlcHbEu1au3f+LfYg1
7IBM4LGaptClsk2LFm+kOPpxq4RQs3pa/gmQr/We0Ufm82YSPZobWqPpc3hZsXc7vvhTGf8B+Ls4
Zja0rsol2yqqS8j9n7MNgyhD0pp4tHkvjWMWQkHya6E/70cFJfSIoqIpIpQiE4xaMTFtkpmAos7+
h/D1LfMI6IBtgcTrT0YMvzBBXrU7XjmKE7tKEIDKzOkZzWWGqjK3EPBHSu0Wh34dWehmLIdnUlas
SXZZ7LwXxEHSG43xNNmC6RAba79R4jTtMyvF3Rt04dCFf2blHEy5I+Rc6cLv9nyPYZdkCVPCqa4m
0j7DAJJxczkKqDW+ivvjCGV13T1grMhO2pGnuCz5I4SYHnjPFraw3Tih36A6GLkFYK27WrtgBHSb
SAkm0+6+qxjNDn9rFtFSWt38EWJ9oK9NlPjT/oiotuPUtcNRPfAgcL8cpQXtEcBz8PrAE7BcmsO4
nUEQwEhB8K23DsjWuPBcn67OROqR5nHsepvfGwIQ/VV5msWuGThy49P1HJeeo1Ez4YyBGTsgndY+
LiNFUiDDOj5yP2jzcF7oqnluyCQoLBdrL2iFWy1ylF4p4BqNHzmIN5ECTRBEaW4wHEAxnmcTT9A0
CHgaUB/oK/U8a06cVvTq3IeYpBofgB00VslrajTAWuAbk7dvookz4RhhxVSbd8Hh2QiEFQeEfRet
6KrG4mPQpbFQ0GSF6U25hRHiMIL4UDeoRI5/jfsllxae4WV3/e610ASG2FqLREBoDM6Ubog4eONW
nI6HB7aiucYcnTuz8y7RxwrxWlU1N+JVajecHntG8LUXlRZHImoFkVDNTiRaeTBkSTa9alzmezHw
lkRD5WYknAZOk3lSRJ1yL8a3fLuqh9ooFCZH1WBX7c6cr2d09X43IW39T2vdnu5U4V1RufYRmD0Z
lVqREtrYXPKPOojETItDUifVJhJVpsaqtEWhW6N5wFsCeuCm58Bt8txd9RSjwcVKdSYw24IFV3YX
LhlZ2BQU/qxtr8ItyaKpvnIQOPXsPfdAsbXUj9xQoJA1qG70j0QZsM9TmEWdGHNrxH0clOW63fc8
P99h4EL3fsLCe6HNwHJXyYYZgtO6YX2XkNHUGFC6ShR9StDR+z6u2M2NmQ7RVd/nmLxKyneLd+RY
kgtGEaSWTZiCUqP2Uve5NOvOsGhO4g1qiJlZvIX3JbqK6aG8jv9CC9KBDiyHlwOp40y4biHxRvj2
2SnU5QsbVgDy5jEXMbfBWRxSMqSXbSDCK57ZqWl5KJksS3Qc4WZNnx89dpzD6Nfs8pZQDSQNd+EJ
OXaLEfKDRbCte5VGCFMQtP4+nQ+yxr+5tuAQlbQL0PoI/2ITrvCPu4cJxZVWLUEpjM5x0XFwS+yM
AkMSp9ZYCx+VNP56iSh+vgf3ALiPIkrpfZs0IPHlmNkbx/PXCMcG/GEpIzkcpCNjX9yDI70DTk/x
xe6+ieUrr9g93qm+9yuW4ANK6G8v/0teKoJnOB7mEU3bkDrb7G+kBIhT3ACdHjlD2d4wet2hmOdy
zPl5Dhr+bNH7dYK+2oov3XlFOhbBvMjIklGeM9Xn4a4ZJVIBLo1/0spe8nUlN6AaKnoY8j3DltoI
6xqpXdKx4yLwwasW8WMKMhhqoJrSN9vvrsV8ItzpXdGzWU/rGeaAub+SVILcHSyBr4+5ZgNydubb
fP5ITKC+bhttTj9Fy8cj+mgbUh5J2DHFtfMLTo9CDSS5yWQpjYlhmI8MbhQ3drAiRAuAbTxdozDV
WfaU6R26Mosb9marMGG+NtIDA0vG4P2NHZcBdVZvnkwz9Pml6wf6j+7Nsh1Ncl4NYEuV1P1PotHs
8qyRuGy5ofxUc7oyETMfb7sOOJkbZQz6QlXxMzQf/Ee+J+0krZrp8zBHBSJBeuGrR7K+nVBc1gdf
X6ziRm12mGs6jd4cYuzvwEqBE1E6kgX2rfV9WDoxbJs6DKbym+6yomH1m9ftrM6J91EPiv4K3EsL
vs/3Vu5fctG36qkVdNm9PH92vULSNn+FDMs7MNbeF2bw1l5/tikzqZkF5Jn3mRvs1vd+ULsP0N2R
quaQCj/dy60s4uDWjMgxumZlIFMcCOrCJolnY5zXKuCUc0NSBCy4f2gql3QYxCOLxV0+W33LetJe
ct4RvKiKoUaWMnTIq6k3eWADq3XlO8kXidP0i/VHZnSVjQdvNe4o1TYqiD5CuKcv9t1NttYd13AU
amn6xwHKIh9hIK1Z12H8ocIPB56iMDklIpzvMUtNmPaXDP2T+8cuFhdoFYMeR0NuAZWDZxG1ONAx
lZsVKv3j4eACvtk3BzHeuUPmpIzdQX3FyPEROp9L6kPmAa9hVfC8t5qaOs7z1vkA/lCBoJmmZz84
/OBOVj2xlIieLdZbxhHxl10bndowUUsQ/PlThlcZ7zSigg2suCBzy+Ga9rdfRGAuruzP49EfZdyM
WDNjAQh7qKROS+TO2DttUCq5plbIuRN5BiVjKV2GU8HSJqSdo3tonfAFyrEfA+ZQXgFw59mKTQZ2
+By0VQ/6EWIGJysSNKY3iLRyWuL4PnBOoxza85M9IKBxULTLP/sjLWYxtwdd2CIfSnJX8ep4R9W6
/j7HtNSs3QoOc1ITkEXKZjWsramdBMzxx/EK+SKzlQrRnC7g+DO6WY9sx+JwlXbrh7saDi6peul+
pQIgSgsLMo622vyFSfjkILV5TGfHcFW0lH+ILq2Gp3rOblD/GjWI4Q0tf9pYagpoGUfBFaAKv5Ux
CuCAeT1Ysiyr3cuCUQJx0GXjJTmHXZOn0c2ysvNj9gQUtvnUfCu8MK0j7Z5J1eWw/tRF+ZFNUxRT
sSnZRMvnethwKkNxkAX0SnXirpyXD3Q8mCsIWoGCv919w1pGOQqB/v60ir7nTr7QzusIU4kPZ3uo
yqbDgOu3b73yhL7l0f7gIJ6YsrBrrW8CltonIgchmEhD8th1dwsIr4cOufAdVFXAw819mKTBRJ58
IXpx+EINxdEqrjNhVjGCvb+zgNc03q5zDWz069ywb+WurH0WoEZzkLlpUER/7tleq/jwhXY/UkwY
dTwwxOuE7hCoQAFF3kV8+hdNUeN09YdznVpBw4Wr6prHVYREXZy/AYa8gayP5HDPrLsK2BcQlPdS
PPZfEBhwwXtgAmwWVoEkznkOJZEmDtRDlBEbkLV/QnrHG+fZ8xsdybYezEMW2iQ5jykTyenD7r/1
h13cPsBpk7jeLkUA3LaXLIVJSCI1yJJ7V7GOFtbv/GpciBlQumtLLcR0iPgJW/KbJtUxic20qLNQ
v2qqAV42k5Va2dWit16yodDH5I/hGoUvBIYrk845hokMadutYCjOpfwWLeYjXFHt4un5BnjVAHWI
RilrnS2KVEK7/WoLEuzlt2iwLEtz2TqwpV9q0kHeBUbsxFYnqYXTeuJLqKN6/oLpXnNzi3qxDJhe
j/36biw446FRk/iyVoBJXK6DOSQuCct51u1nCU6AWWujpleE/wVRcb7o1QpKM6yoMmZvdjIbQk/D
RP5rpbuGXeOlQMiw8qxazADrQAugUpe2LwOTF5zRCswSw6xyRt5K9RIP++4BGNwZebTxYLE1hosy
f+jg7E0ym/q9E3xAV5n3TtnkICs26FJPLcfUAgxe+wQqlxjZ0+NFQfgq9ruqPIkQ7Osj/9luwScu
EaSAuLe1VLsHrvx4QM1FXTH7/5SWV5UfFMKhTvLbXYIrcZGNA3X5sqLFulZ6a0iu3bzAyjXLpzuY
ZKYa/XiXRIEcLMuSsj5uoyFY4LKwiqWCkK6pFQcxj4lznnozj4SQ192LHQUpq8CBP6p9jGd1fE92
MiBt5PFvQ6LjlCLD2eZ/A8UjYA2qjV4gA7+hCZq9AfI1RCGiVTxTZ9Yh6SnQ3hZxvsDa8LcnSasu
1yiYuRXFgSAObs6zkwRFKMdWtNnpD9qLgECfV6T/JqJMlTmf08vyxPzpH1B6/abGoDF13yiQFozg
9dYir3neQOY3Ck6HMHa+zeIgdQ9Xj/6VanyeikWH1R2E7G9I2gOdpYdrQS/5JLW/9q5e5JQnlR57
AzqYKKbzPJwCbbvJpGPnpFlsq0+CZTybJE6whSxtSV30bWVfq6+O/YxyEpAwJAbyghWOYQcH4c3H
w4QD5GP/o3f8zXLUy2pMgzvhDbuSlYB7V7o/RH1TXINlLNebXK+eEPbnx748xfw7TpkxGakptYir
XzdojdvZhH5xXoY+HR3jmob0C8jOJyR4oSzBQiAQGriI4SoEq/mhpTesZYxrtaJwV4NKc6157xd9
5imKcJXzxWdohCpvpFG0I0LRxYrRWhiw2iK0dZosq9nkF8+6+QN8K9hYrltK4bZCjIwXQhXTcf8j
+Dmgx4XOD/Y/0Ocm5ZRMihWI0GRxaIEIpQN+1zYKyNBF337nAu4KIdvtMctFztsBga0DAewX71kl
vhSfR6Sea6YqwHZpavuAsuAlsSXkUaQxhzVjn4LWymaBQWrNgSZujZai76i0qhVphaQ8kKtZv+ac
IcLX9C/RWIM0pao2ky1ijgBNFhcDNgjsBt4qd7KfWSp+EyqkELQWdmvAnzmOnKDakkoFnj0m1W+X
nPxpLxiw/h1wNMuv40FhFdj3adg4CBgKqoSE8MzkR4irqvshj8zCUCJjP1xTCC2WLNAvY3Y/F+nE
2vw/95CQoqiuXMobIgK6yWAHk/U2qdK7yzcFHiX/Vlup9BhWDvX5cvYNumE0YaxySBw9TsniK9Jk
FhEaNXfuzG5Vfj1XnkcV0fmJVfnLcNldK6087pJ86bm3ivJ6v5rgku2CcAzrYph5lF7F4ppxWFpF
zmNqLsELXnSWsUnHqErbIlFRqKbF1Xj2Y6QH1ODiiFSa07XY/qvCGem6GV+OqtrJ6IpZVG4l9+aU
W/DHL9VS1Iw1iAwk6UmkStjM8oUSj+aAHpgiL/4dBHwYVOqluiypt5NJq2fvqzqLw7POATOw62u7
gFHSfH8lGRJJ3+v86ifPCnyCtd1e2NYwoZGS3e0JO7G3WfIGqfhSeygYDir6bmkCVpo8fyeWWvys
YAKEwSsLUlALDEn8I2l9o/PF0y8oksqkkou0Q2VMO9QeeBHsQpZtgpPlxpvair5jAwkh7CBuBL+r
ZACNBsesuRPrCuxbr5Tx1n0M0Qs7xtUqtAQMlpiEoVayDAs8VL0huYCgJBVSYlDWz1KIxlFdPDUP
ufDK4ENMofnk10c3PXrFf09JxX7+qZlwTRUQZIq/YI5KxWjM06JBSu1nx+wsbbrBHs3A/50JTzML
lGYK9H/Yh3YE3tvggTVIckY7PKgAAiQubjTVxarjlOJlgx0/CkAtQo+Lwf8l2L8ICG2Bol+NBmfN
Ne6dx4BnLvBRACZmdGcEwM46TkS43MWZHeJDf/oe8hW25N9nBZawRMd7+iXy+fjIiZZCW5J5Avii
Fhyc3HQ9VxWdkFjiZXH8PcR+BykZienbtLqHijufyQQk6HiSD2E8l/yIrMOR2rB46Bzxz1+Q/mQC
q0mQDPcEDIqFIibuGOUun3d4815YDS+Ao0F1czpkfoEHUStp6h4AZmSIt+IAhVQtpR39kznvuUzF
zDl16XaVNULeWbnd7UGhQQN5rvDNbuNJ8HBPNZjBNPvrFKLkcLNZio6fJNIuRDTzKQnFDaXOkFer
nK0trE8vOCBjPXQtffta3OwO7TNKxJtSH5yeb69+B0c0Lz6TDrpP6Srddg3uk7LTLvn5QyBdR/yj
FPKRAWJTW6luW4Drf9uVxfgmpy8pULV3kOH+IWSpkw3Bh3bT59WmLbutsFOA8fY7uHUElZQUs6aR
DdB/oVhBbJy/y+6rbxPYyVG3Z1dfGl8iIsXqBm6781DfXNp4bOnbqmKt8QZT709FIvf4I9lLzwPB
4B3vrLSF5D+x+jEEDjUyc6NdBjnM18YiN+BEgp/MxnpChFCvzp26s3UEDhoNLvG1uPoMrsWW7wHg
n4OI72G2B909UEtJkTWMyEBvBNOH7DdCIq2I/K8GlziQ7IC47LrmsRCOCOv7d53mqa48dZ16PiCd
i8vslWBe0iklN84SPv035sVlhwH3y6j3F59LPBwYm/q0UVxF6zbcgH99PALYtd1QGr2faGXhIV4l
OSEIS6TvND0+Er+fsS9fgQ9VFDOugk9zVvzQ3W3FNQjGRU7E+OhdjL2vzj1eDrnD2BUUDBJZyTQ4
gcEIOhr6/yvJs30wTq4LXE0DIIaKra4Ejsm9pJZiZxq6pNlz4DIviBAgKoqzL1WqqQOJIYMohQVh
lcl3/z90R8QvcyJ1offviP9C9T6KGSfIPj8Q+J2nP1pzOXeVGObHcC8h0sIQzhF7cAGSey7JHWou
vZIudzbf+LPT+QklaRNg+4VYxCoKqKXeXL7w++Q3rZLRt2kKgEKs0UUtZoCKD1GqweOzcJWkBGhC
vBxF1XT23/nnwmiRJU7uYEXZBpHhnW5eAis+kCdMXDJqmbXAjy7zV7AkR3zElQe1ZbMFejvp2olO
4/JszfD8PI4gyz6W4ybkxGFjVTPkamWYP8iy5iP06GLZiiOIzFXwtml+op10aAxE2y+eOm/FMn0+
28i7c5K+q62wVbLvWbH24UcEi7NcC0+vut21aM/3cE2UH5fgAWMMwNwgb9nCgPblAG8xW2m8/pSm
mDUGbHo2I6XWcbievGrUMLQLG6N70qngfycQZxK7TkbvQVnkXxxD3sCWiKlgps4B4/fdSO3bJq1Y
PtJIU3oKZb1NOVbuQrmkw7OHoE9Rezlh1ddxLxwQ+SPaI5JE+AnO3W3nUqN10/QrTis9BQ49UHZB
Zjufiv60K8zqFJyEfNlXNr7CRuVzNo6XsxHTiGbSBq3Sd17KPGtTZopqB7eBNe+COyhOAJkK+rgv
7FVppt7w/Cg9e4PUb4CWCVltcn0DwSXXsQh+uF6G+Ol4xe+Ki/9/Dw2hfduxHKSVof3koNvyEQH1
ZpZ8sDCfswNfT2aNtk1esFxPXtuk9vt145WMB0LNh1X7WoQeNjnULQdazXB68dESGIKmh7Q1ncla
qiT5HagtVINQRJ7dBG4qPww4cdw3D25+3YPTJxu59AFXKg3GtDubGYx2EB468DjdL5Y0JweNVHsn
J5YjKsiHUry3pdhxi9O0oGOW4IUzz8cyXVN9IRQ+GAO1DjoUh5RJF2CeBIF/O2kXm48bdbP4h4j/
wBsTkfj7VeRGucrJU7BDgls9HuID4nC/ykzWfo20FCarT5SyAvA/8kwK1637nN2hbCM1iIs+uYvU
O4i+7RRgiK5qz+aav3AaAXwvcJFy4xAnKI9HISstkRraSl9dKBzbhp5dxKIzRR2aGGBdMUZVtyEp
21ozpBosB57xOPSb2VWosOJe4FNXCxRrz1unPLzvfmbMHYhX6dC8KObSjcSj/hC8xviVkohSC0Ye
TCQDSV8gHrIfjuPFfnhA0TvUXeLW6O0e7OdsOHDa71XLrsc2XfzkxpqAspO1xixc6rS4ZIZpStaR
dnYj+mXrKqVthN/+ud4r8bTjWu5f1Up1DMs9dQXeKJUjSGSfV8Dwri4z4E8UNF53RFG5uD77Sdoe
9RCQh5WdejajLh80SyPtMo6b0Q6SKSizniKHHSrrJ9wvdkVZsnguja4Q6KfsD20yrCvcgl39VS+7
P+ii1EtPPZzHTq1F86/ckt5iipdarE+z0FDMSr1kmUg2hxod+ObIZtpOfJ1d20oF48cV/iz7imn+
E+GGMfkDgalH3667kE/NdDwrIfRsR8Suxis+Tlpxi5+eTPLcrWF85L6yLD6VKQu28w447OV8vt4D
StoymCRqzb5djBZOTWzYMWdPp/csEj8NWFPJ5ctBUVYUEY5nQHbFghtdOZ/RU42kguc7MNN059jk
r4iMSQeKt7u8eKCMDHAlzsSgC/dtxHFgsb3o1aRTAxrrE8LP6b6DZPaCwvwS0mpx6EVBHs7pYsor
+DYauUWjHfxR2IgiLzjIMwOrvsOY2WyiqBUdiWyhOFmj4gLV84z2aIF8bicQET2sc2YYus06vPjd
M/seChwTHVMMuVlr66zruQ1/j5ns64N5FWpx5W9++2fHk35iYUiIXm8nrr7DI3H9K32Obpk+w7/o
7DhuZE/38ogAgmn2zy8DhPKSJGR4Hp426RMK3LRKq0VgzHgAJEbXBB48uwS/VU8rhF7xvf40y0T8
YSoAP/sc6sZe0rHumz4oYceGDVItuMuxZ+WehsxqzouBvey1pNxYSeJDVkwuIiuEwPW2TegTWkhl
hgnx0jlnxKmXagy/1AGLnY08T/Fhyz75pUWo2wCfS3tjzKgd22MS3NramqR+0I4RobNjYXJOaYMD
/ok6n+Opq4/ySWBmebiDhP11enRnTb48vXo6/LIIg9/UntHVClvRZrw9tnuaI9GpI//imMzcwxbl
75JcmC9XAMW3Lp3YIVz2l1wV8e2G6sVR1s9jnaczKMIh4W35ZOl51PdxrZuIf3NiPMgZ5NcRdBkd
mhci/MgU7nxq+v4Tr5Rav3DbYXp5SOz0hUa7D4g0CYk2mU+I4jFYinAU69ryPOl8iPG1Rkq+lF/l
v+gR6ySUsqozOIzjIOAPDTqIdZb4QIVBJ7vZhtK58cSbgfNeglblSQkPEQ6Rsuwv52bkDN6u+P+S
aHkRJBa+ThHX0u5iaB7cnPcnLm3cETXgOWDWP3Mk5PVQW76olSeYJMFNMJzg3/uafgXsTPDNOHl9
yjpaFKyneDjrQqEBv3dD0dg1aZ1CzHEv1gzG4uhIm/jZRQ1pRIQCDAL2OYOiE2vVs1n+jV0AZstp
MyxU+QszZGl6nXMPtPXIVDXaXmDZ1co+TLMBgyOqpkDhIXXog4FlI9OpPDtcjtFdsZWQMv2j35wA
nv4wgnVfUIPvJcgxvhBqvp4yqSoz1JyNGqnSO0QKf0AcjfXhERDQwhUYbep08rYHL/BORrFGQ3YF
J55ZFr0qVb8FvxyTdyVZLE6YNpoVHGKbTiHzMDxrG5o4SbrGUPpRxmnNF1A9TqfJGBWhW7T1y9sd
fk3kWjiXO2zAicxIqx8URG4VlUgf5AV7wc5JlozUj36chAd6w9be1SrJLksJnofngenn2llugwR4
zbSCQSH1+qoPDUgOXOlJcRHKVLmmeuNjhqcMBtS2ywQwvud/vfbtxPIZU3Gl6USuQO5HBb11+pwh
GbBKiOeAhW5PgeUrlXZj+WOeDghApanpDeE68YsCu/vR9OAGtMT4PktVNQGNEfKa3+WFuduupTJJ
5PwRY8Ga6vmdew4Scx7yrMGLQsO+MryzLUCD/HN8DPY5hCDlgJOE2qKxGe3ZzecPWdfe0kt9lPBx
fg8XMH+lylEZRXdXt6Uwb6xZn3xJ7nQtTFohTD1U7Jb0ZLA52b7oY0E32fAeg1ihpDE2k21pom1h
qx+AI8/OXkHxrxCDDQQekv3g6cqxxvLeDkTSQlvFjkm1VUL9rSaM/w9o/dUaDeCH3bLrAfSi+o4I
ZWdeAsFeKXV6bp000b9N3LhzHnZWZEy1Nq7NGp5KUcfl6b5q7BgAWjzFxU9P/9jzIwzDeoVYSE5n
nu9XL5v0VeSlveQyS8/HMOENCUYfk3FsneVn+D7EyiwPqlall0K0/nmwr8p1o27HNo6GpKbe8s1f
gHuSZbi4BoXwGLVAFFKv4Hl5J5JEKMRF9R374J5nf7P2xlq/VmnJJ0w8+aV+fnL8MEoxxgGJ8hjz
b/6L1Q9wWmawbIOUhnmORiP2ZHzSO7v6k5pZzL7ZmCz4qpPSr+wtIN1ooc5NFwLWMIlNxqx/O4kf
FeqWE2mXcjVUJ7b7L0xZnqez2kq9iPCeqUG9hr7L6XzGa6ztRqNX6lxJ8DzUAf/Txl8PE/f9II5B
OsyM1MKP68A/j4olg/oLZHLokvCP27jqCUl/TE5HPHEenkTAtZhb40tfkhhgPs8JZBCS/OEKZ5If
bDOsBJX9KYa2pBfmNW3UrJj/R7h/ymd5snM75ebFVvEWHLMN+hVT3HS3fmCEmw1bc95+CGESCgRx
q6nEj6Bs+CeBnImOYUo68LdDCK2us+StIzVFoPjT3kWwtlBgStVfsLS4sVrKUDJK0Xx4NZ7xXGgO
1baJ8KtXxK7wpvtV8AKMTdDWaagYrBe8v3Cx89ut55fvOdpVZ2v24hGeBP5B7zJgIvR/2Zr9OUMw
inajNCPfPK7iD3nRdbjakX743Ol/IqcN3bF83dnSlOjmL7CaTBsGMLS6ztqyQy2QS561ltGl6tPa
UOMrKAzchZar9Fs5abjRyXvavk1hfzdYBSN9NW9uu2NpyIr6zWso4UmpZzQNkVyNxurtBnDgNRIh
Ii87t+HgkMJZKl3DHh6cLib8cIbrtKQfjbOoho3phRohtODlw57j8zUBGcwui/t6G6TEL/trf4gX
SJK2aSmvYbBCXvJpwMjRnq/EJebMuuXSNLldLaC/lpaqKpK83ddsX4qeAIi5TGO9arj5N05Irc1A
w4u41qxpegrcibyy7328pPArjEjQQzr5/aF2SzQ5DxIqzRCB2kYVjf2oEwLwTqV9dczo5SrvX9lz
r+I/DBXEOhQAiCF+y5gna/HEekxJ9vdq0NI3gv9u1EmVwkI5rW2uqTqlUx/tPZb46u4gx37Ul5oj
VJH9UjSSaUBc0zcP+hGlDGQ9dn7/LqQqEseZJzExz+8ATfJUxRwRyUgrk0IfmJD0TOEIqExhuWu7
UTuqXX5xbzC0qJmU0L2ECQMBnPDgRyJsbLynUXH8+DwXR3cTewGtKgpVbZVY8e9gcb3IHZlw5WtZ
xPMoKsoCdI8bkPPkz0NzFNHCNmL5TvPRJ5/NtnMtqrs5ROywjmRpjLQ+2NC1UM/bDcf5iIRavqWI
P6gkM4xpMFqQjvsxRYZl9SePHJuG6upx7SU3jU4ZCrc5sHrbLaL0QkB6VKvMpbEP17ygzHEtXODF
dOfjrQTCLxaPUKLv1aLy5Z6aERo4fwEnT2R8Hpbp/a/zd3JmZUeku/aJjlmJeeHit1ubsljnn70e
PK/hgmyxBoUHQ7DZlmFgQWmy+c/J4xpusMV7QkLnowE6B+1bTABTshzUV9NHONZNeQu2YQOqnyut
y4xm/CKwTZVoXaRr/UlZdKXqu3DWzoKzKKOp+dUk6d7eLpFuE9MZydhWk1cdImXV74Ixwx9WqGHA
ky9XVE4+W5uyubB39zUzArdJXij1of+YGg6vlmGIFlQxvxc5H0PbsGxD++18QZ8D6Fd+T7VFAfhn
6a08BXpy7Qhr2R3KPbahwOhrwYxAFwShAobjuLbXDewFjF+qVQOps3qWNTqT7n98ocpVSjSzqEOq
4eO8qcRAiZJLxHdeOcui3gnlH71cfSzAhyKU8IrJO1qFQeUHlx0f24HxCr53XlJIot8fQFHk3+Ga
phj4PrKtJAgJ6+NfWWdj01YXnb5ZLegKpyjLJjIb5P6nJ8/XC+LuQa5SUCpwYvmlBJ41iPWgEKnl
OxAE9oTmqTvPvnyL6rBtEKhEetvC1mIZhYVTtUPBQxeyMDHqHmAJTdL5/SU3Hp8chbiuI0QUCFKk
yrsCe6oYCIA9j+8k02ge+TKpC4zfrCyWhOguxehclXrhNF/KIV3biXYn4omo3ehtBMktpFVSxqtA
kWtiNcGCN1gLmsAq6AtbFiHztE6y5yVaXffwti2Sg9hZQ/6S+752YK8DQuZ7jGYVFGos8YRHJT2t
NoJo6zvx+tEmYgVYJAHpuYumq9upFsXbT19CQnNW3j1xvdUxbsz9csdBAcZLe5yooLOTJh//7kpR
0tzi0AYij9bKbknEUtSLh/lVJQgPlOlNmHnxZwMs50bsJdoBUO0HfzkNXWWOSfsREdUQaAhB+B6b
t+5/e9U3j4Vlletoz8tMeQKVIAmb4uCnY9edXar/gzrAQ11QGF0EBcbrfUvToY0pu7XH3TXr91k0
pIhqFQq6w/LfU8eExEAX99toJhLwzf5AQWqX1Y61EGmjrAMGxw4ablbLMV83TtZS6tro4Bh1cCSb
ixWmUK0f6eIsyko2OpYF/YH2YKcKu3RWUQXVI1Ih7qxV8vRUYbqNGVJWVkvX8FbYuPKbQOhNo+aB
7fg0mHLs/TRbBAmz4KHSXwiQ8x7vi7ltscuTBNGPmn+xWU4vYhRX5xq1AaOGfLWxDUHp8/MwOcZm
f6zw+qy8LYLoumTZoz3UNIUoCmApJCiARuOAKMHd3Uq2Ht1eNKXdfrtgDHVc14DWilnLsqrXzax2
bzekvX1qplnuq9E1+wXQpM+CIK7nkhElWQzHKE5cCBkBdpXRBRo8IWTX2JEzKVhwmal3g5dr52NH
PcJ54Hnl4Bw+aFKaal5dW4+oDwyAivDCEFdbTzTihDXzs8quS5aczz3hGTJ7vHfT7x4J60wyeSg9
GBSGkHvjjlhEPyzm4Q3jmsZrahNKQM4XQ5xEs9AzVP/vCgqbzst+BcuRlwl/jzoMdWfp8Jj062/m
2M9f4ipQgos+xOJm+ijIomibcnIrQgSoXIE+PugBApEw0b+X6kfamQBvg/l4eZLKc1n4c5068KG4
5uFNhTD7IHe6JDdeDWOz8mcu3tYiq8MYQC/yfl6K2Akmsw7c/WGoyoJh5SsWBbaFQTp6LRrvGLel
GB0ntRDDa4nG8GoocCAAlbqMzlPwSI7GLwpfPW3/sX5B7BGrGsn+CZsppgv7f3JcnqdE4+yDejxz
YysxYgEmxWPw5lRzxEttxUDKW/tDFmMUEKRc6Dc9l7VfSq55spfZXJdO6t35w/7SbsxRIVAIeHgS
1RN/3YoUAKwy27y0Mg6h/6xlRdaOo7ueT5IansP2rwO5GAB2fAlCohuco4N5LLb+CHH+cl2yWalW
7qKHLs38ZXf3hN6UbXJvtDTu8C4yqOaHTuzPPW7sMaQo3jTuilyk2qMOWe8tU9VmtN3wniaVczX9
KjFgDyoHJ52rDCgVlGTb3QMVcHiQBdmeJiinZGDffH13JDVDLZ/FfluvPlXMR/XgjKW541VOH0nm
OSPvS9F+g3u/N/3bzfqdzdrOLEQHCA4ILMU6pfLpcjxP0oYySUyKGmLIMCKj/g4yVP9dr+ukz0am
VDLVaGUEbqK6fR8TdGbZ7dcK/Ebg1qZRaeRZSjAqT8alWx9SOOjOcI9mR8CEQy27IvUDEvHsClqV
HjNhl8mtR1xHNIHwUpnD7qs22+Ouvnhj0EGdaswQLkDyShGCUfRYZFM00RbX/VfItltPOpW/VMCl
jC7Xs5jBtrX93ym5URc+bL48GthAr/Uk6BqeYibr4HSR8yg3/CZ9/MCqma80gKKQBQtJQQv0OOl+
mWTq8S8NMX1bFonQqv7QeRbVQXlWij4gAZ0nhXDqvcwY0k2aLX2YiDdK559Qu5Oc9+kIJ0AWX0Fy
ygrPNs7XZG86JdmyMrTdsiwkM/RwDE8O12fZkCDPcImHCixQoNJe3AqKwlGje0t/hjP44msPtr60
T4b3tksHsOcQve7Cg3YwK7Y6WcQt0W1UcDGa/GVizypeVaONrvA+htXWzCGUXrkQYNvFxOGFk2fV
XWs24DYnVKaaYnsJaOnzBKegr/I7bw916rbsI4qY91lcjge9GeONM4pxvxm1xx/p/FrCieYC27sO
aXSectwGaEbI4iI6xvw9RIz+KJ8k6mpfnq4sm8CZjUS2k3UgERFLCp7BUUELyQaSpPoOjsQZc24O
PatcKvTKkSeczN7J6Bo/KCYavC8r8tD4vbRr0FyYkyHPHXJ5j4YAK4cOZDRttl6atcagLjffL3p0
BDkC3YAmF+Nh7p24KY7DcaXFw8w+rst36GtAuH9Yoqppr91WP4vV2V0snvRuUZinhrt5apwkFI5p
r9+unK0DeQigRsSW1lI9OZ8ON/oN4VA6ilj1HvwnfOHhXFXN+imQoYFJghhLRiUBi7lVdlEoFjcH
4vzLZb1HCkBHM3kdZ41i8bLjnWVKGzvHbsC+X8jBsQBA2T1+hDjcPrkRDQjSoe5nSpBnJS2/6rzj
Ou0kplXBXxtUQ3ltOo3CY0C5ssSJ2lzHb0rIjdtkJsG1aqWbXflqAHKmYQN2/kTujHXzC/40FUDZ
52cdUILxuXHGUPHoQ0jYVi2xoMppk/Uz/eg0ZUaqRNGriws4XXb8PV78ulU96C9Qe89ntYb15a92
Ll09193+fLhQGZ/8MW/MakQiccbj5ABK6Auy1qYX8xdSl2G0gaDYFyv7sibMMR/WxWsZRRzZdN6Z
gCAlbrkp4gBoP210hroR/NskDPuZ2vjXJ64JPirh/u7jNyznke3SYPbXBr0nH+zQfOBrQDVpg4kg
W9PckqOzWZUkhaAa3pohdvQ5PsiEy9S+kArLt1jqSETXyWFEu5+bQYsh5XseJsdENjryK6Qwuba8
amQe1OSE6Sg/A9RMtzbP9lH0GS/JU2m2ZkdvWhSs9nMQVxmxh83InqQD1AOXY3YlTxmcsN52Btxp
OmpKAZpM6L2NXn1HYPl3fzKtuj6x9Wv3eAFxZVDeB+eGGO235wY1Uo+iVl8DHUz5Pfz+klSzq8/d
DIj3g/mnullfXOfw/xWLPTd6n2AalQ5xsOeKhVkVhTilowAjBCyRTeiPL/wOjcg5VcOu4t1roayk
5am1UOPQkyD67f8UEv4f8NIX28bI5tHMnbdO9I3SLpRsOkOOPIG/3P9N2O2lI5yNZKngur9xb8Mb
A5Y3iKV2onAO1hlN3jbtZGxLWDSfE/8W8w/NFK+Biqyrv4lgaYbn+It0yY6XBr3UCxkKQYZdAKD6
kVuYUUgzvhx/WSFgvGdqYS2+5yM3l62C1cl3YPFbyN3VUnbGljFa1HxFEJ4Y6sQ0T5FrJCkAECQi
2pW9i8QsYU0BVy0HqyV6cHlSjEZcQenfkggpKAzrl3szkl8760nhCmbhNjFiLtkiSiMxBW1K+L/m
AKRIS3jWXsD8Ka3GugI1+SK0Fi98E7MzK0BuIiKeE5ZcqKPW5ig2cZB+5IU41OFC+ljGXwZNIfUr
8/jIBCVN/mUD93OLOkl5vXyLdbHXD7lmzuc67uXRSx4IKzW5s8Lq5sT47fO+4qe3zNNACikjoO46
jt1Li+gX/bfH6gWD0XaZy1grmrVU3bdUbWJg0/fzkQDS98I7tn2szH7YO/xFuSW/a0yBfIpRwcj2
t3WY99BDrNS0SC9FeRCxydX51bOgWJGgxS7tAZIDKDG/Xcr5grpfLo9hGdShfR6PNVVtFnigr0lg
fGAg5OubUSyxBueXGat8uBbD0q86AvdDeDrYCvSP5gKgIRec84Ga0ocSxlfhJ2cs9CJ5BoSl0Wqe
+Zej1JJ0MMvKCV5X/ALnv2xiyHwddOfEFMSzWIcmXNpAno0fwbpBr6S5U6ANiymSGvYcWVrAaJN/
Q2RIKi75TLrGvgEXBvRsa/pwTCzaxFI2yx08xSXJ29Q/n1iCPZjA0ICKmOTQtlRErECeo9HbG86L
2kCMoUZd7ShhnqKV2bRs8mOP2Ju05wvXVvX8m1agAq3S2SC9V791x3Il7RMF7LqCQcqSJuGFXPvF
jldyD1zlj3+3qdr+0mr72SDjHX3w2g/pDRpS7FOVDbQnNoLQlAsXXUV5zoP6kTL9rBK2+nqy6zTD
OymdF0njP8LICveuRiwGbFhCP644AJTv999ttxsqwXrO174UBgLLgNdqPiG5rZAn8Hx2v0cZEhmj
wbAxvZGKReAiO42rHLXaIjdcpp+ODglDTceIMNyTSi/BnS9QOYor6aiAGrWfNtfZn3tNrRUpubS+
fK7zlSFvKYs5HwUpSPLDAJH40N2gBQdFDxtJfr2ynnBC05HRFsWyvOWJqxdouLmsCooaYgPLnIl/
V0oriWABCacnZ9gI7SYC2y1OalMYU/4OrD3izmiJHnjrLF2nB7XBxskOesGHnYJqa6akqMTwMElf
l7DRr8oIbuYFHy574LpadCDg8bN/rxlM/zSSV+BcF1pZQV8xeu44wFq3fFG+a/YCLfczhQ4iTaY7
yYFzSPctC98NlIDYTPiqqI8c6eekSUBJNAk4sZ3HJ6PBjB5sPt00gWXbSqS3zrUR0+hUMh5piYOe
iC8wuHuC0D5UXJTvCmavkB7FGrBmnb+PBbVKllIPJsbD/IzL1/2eimUjRzZKiH9Kc7di9lksIPY9
1Em9tWx7hGv91tKhMwQX6oY8uqIADbe/exwyJLWwsROwVHNybd71mp4W3MD2InHTn7WNDAJnEx02
QWcdmHXo1OzRBLVft6cQ+vUocsH2aeB8AObSaQ5LHQD4+fwWdBJUJ6YzkIRD4EKASTldhvBtnFgV
vRd8u6OYH7wCj3Yuc1dmARox/13GLfWjBabFxj/YPfnfYSK842YNPib3JnjOYQgxXvr3f6dHA35U
T6K6asezWRCcxRagkNpeL4B/28eNEyVJFuUc4CscVl8zARtC/iCAtraRJUZI6SgvzNsFDkZ5XuZd
s1zWy7txpYh6y86yPCcEosAIIqc1c4z9UtwAqa0jezAxJ2rLwMn3I1WoylPwPJ3OTivsJldgewPY
KHfd9JI9dr/+T1O5Dvp5iz7QYa1YxU7TT11/0O8Vb7Rt453LU6dAr/9W+XSnZYH96etHR+PnvYq/
iADQO3TndUYZQZyZP6Mfxq3XbAsscO+JBs4mgqmxQQCqUpEM/KdFT6JYz9ywpNz7dmfilAXO0Gv5
6fcC8LqJQsBSClvCusu7JyYkHTmd4fpDIH3bHgm1XgdiQ1KFvHWaznTArdY8jQ0iA+Gc5Jjmgjh0
FUQnF2lfpXiy2GYC9pWc0bDy7llP59lZvthfk6/HFTGw7L18yMXfAC8JsNxFfI9VApJqLjr1e4TP
obN4jv+kgFh9cZCtaQB9BAtXpiwr8kNkOtm/874Kj3SxcupB1YYC4LB1nfkoRMeb7CSCGLZFGqSD
MFuYCKzgrNZzj4K2zCHVcz4xjkua5tQQJLslo01etuMmJvKcj+XsgsJaF8YDE4jt/F6Ivd5I/Idt
sQvCgvXzu5rHqdSg5ZIRdVRb7A4fUajfpinU/IkJAaD41EACWxDWI9yKbUgtHjttmMIZsVzQWt0p
Z0JVdekGMuSgjX7SjAvYGdAzxfHLSlpUHQCYWOyv5aCa9OsrEQeXVVoJTHE3ow==
`protect end_protected
